* File: ROM_TEST6.pex.spi
* Created: Mon Jan 16 14:53:16 2023
* Program "Calibre xRC"
* Version "v2016.4_15.11"
* 
.include "ROM_TEST6.pex.spi.pex"
.subckt FINAL_TEST4  VSS VDD CLK DOUT<0> DOUT<1> A<9> A<8> A<7> A<3> A<4> A<5>
+ A<6> A<2> A<1> A<0> VREF
* 
* VREF	VREF
* A<0>	A<0>
* A<1>	A<1>
* A<2>	A<2>
* A<6>	A<6>
* A<5>	A<5>
* A<4>	A<4>
* A<3>	A<3>
* A<7>	A<7>
* A<8>	A<8>
* A<9>	A<9>
* DOUT<1>	DOUT<1>
* DOUT<0>	DOUT<0>
* CLK	CLK
* VDD	VDD
* GND	GND
mXI42/XI519/XI72/XI21/MM5 N_XI42/XI519/NET114_XI42/XI519/XI72/XI21/MM5_d
+ N_NET127_XI42/XI519/XI72/XI21/MM5_g N_VSS_XI42/XI519/XI72/XI21/MM5_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13
+ AS=2.397e-13 PD=7.2e-07 PS=1.49e-06
mXI42/XI519/XI73/XI21/MM5 N_XI42/XI519/NET36_XI42/XI519/XI73/XI21/MM5_d
+ N_NET141_XI42/XI519/XI73/XI21/MM5_g N_VSS_XI42/XI519/XI73/XI21/MM5_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13
+ AS=2.397e-13 PD=7.2e-07 PS=1.49e-06
mXI48/XI66/MM4 N_XI48/XI66/NET52_XI48/XI66/MM4_d N_NET90_XI48/XI66/MM4_g
+ N_A<9>_XI48/XI66/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI48/XI66/MM5 N_XI48/XI66/NET48_XI48/XI66/MM5_d N_CLK_XI48/XI66/MM5_g
+ N_XI48/XI66/NET52_XI48/XI66/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI48/XI65/MM4 N_XI48/XI65/NET52_XI48/XI65/MM4_d N_NET90_XI48/XI65/MM4_g
+ N_A<8>_XI48/XI65/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI48/XI65/MM5 N_XI48/XI65/NET48_XI48/XI65/MM5_d N_CLK_XI48/XI65/MM5_g
+ N_XI48/XI65/NET52_XI48/XI65/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI48/XI64/MM4 N_XI48/XI64/NET52_XI48/XI64/MM4_d N_NET90_XI48/XI64/MM4_g
+ N_A<7>_XI48/XI64/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI48/XI64/MM5 N_XI48/XI64/NET48_XI48/XI64/MM5_d N_CLK_XI48/XI64/MM5_g
+ N_XI48/XI64/NET52_XI48/XI64/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI48/XI60/MM5 N_XI48/XI60/NET48_XI48/XI60/MM5_d N_CLK_XI48/XI60/MM5_g
+ N_XI48/XI60/NET52_XI48/XI60/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI48/XI60/MM4 N_XI48/XI60/NET52_XI48/XI60/MM4_d N_NET90_XI48/XI60/MM4_g
+ N_A<3>_XI48/XI60/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI48/XI61/MM4 N_XI48/XI61/NET52_XI48/XI61/MM4_d N_NET90_XI48/XI61/MM4_g
+ N_A<4>_XI48/XI61/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI48/XI61/MM5 N_XI48/XI61/NET48_XI48/XI61/MM5_d N_CLK_XI48/XI61/MM5_g
+ N_XI48/XI61/NET52_XI48/XI61/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI48/XI62/MM5 N_XI48/XI62/NET48_XI48/XI62/MM5_d N_CLK_XI48/XI62/MM5_g
+ N_XI48/XI62/NET52_XI48/XI62/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI48/XI62/MM4 N_XI48/XI62/NET52_XI48/XI62/MM4_d N_NET90_XI48/XI62/MM4_g
+ N_A<5>_XI48/XI62/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI48/XI63/MM4 N_XI48/XI63/NET52_XI48/XI63/MM4_d N_NET90_XI48/XI63/MM4_g
+ N_A<6>_XI48/XI63/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI48/XI63/MM5 N_XI48/XI63/NET48_XI48/XI63/MM5_d N_CLK_XI48/XI63/MM5_g
+ N_XI48/XI63/NET52_XI48/XI63/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI32/XI9/MM4 N_XI32/XI9/NET52_XI32/XI9/MM4_d N_NET90_XI32/XI9/MM4_g
+ N_A<2>_XI32/XI9/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI32/XI9/MM5 N_XI32/XI9/NET48_XI32/XI9/MM5_d N_CLK_XI32/XI9/MM5_g
+ N_XI32/XI9/NET52_XI32/XI9/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI32/XI8/MM4 N_XI32/XI8/NET52_XI32/XI8/MM4_d N_NET90_XI32/XI8/MM4_g
+ N_A<1>_XI32/XI8/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI32/XI8/MM5 N_XI32/XI8/NET48_XI32/XI8/MM5_d N_CLK_XI32/XI8/MM5_g
+ N_XI32/XI8/NET52_XI32/XI8/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI32/XI7/MM4 N_XI32/XI7/NET52_XI32/XI7/MM4_d N_NET90_XI32/XI7/MM4_g
+ N_A<0>_XI32/XI7/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI32/XI7/MM5 N_XI32/XI7/NET48_XI32/XI7/MM5_d N_CLK_XI32/XI7/MM5_g
+ N_XI32/XI7/NET52_XI32/XI7/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI42/XI519/XI72/XI21/MM4 N_XI42/XI519/NET114_XI42/XI519/XI72/XI21/MM4_d
+ N_NET129_XI42/XI519/XI72/XI21/MM4_g N_VSS_XI42/XI519/XI72/XI21/MM4_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13
+ AS=2.397e-13 PD=7.2e-07 PS=1.49e-06
mXI42/XI519/XI73/XI21/MM4 N_XI42/XI519/NET36_XI42/XI519/XI73/XI21/MM4_d
+ N_NET143_XI42/XI519/XI73/XI21/MM4_g N_VSS_XI42/XI519/XI73/XI21/MM4_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13
+ AS=2.397e-13 PD=7.2e-07 PS=1.49e-06
mXI48/XI66/XI5/MM1 N_XI48/XI66/NET21_XI48/XI66/XI5/MM1_d
+ N_XI48/XI66/NET52_XI48/XI66/XI5/MM1_g N_VSS_XI48/XI66/XI5/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI48/XI66/XI6/MM1 N_XI48/XI66/NET48_XI48/XI66/XI6/MM1_d
+ N_XI48/XI66/NET21_XI48/XI66/XI6/MM1_g N_VSS_XI48/XI66/XI6/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI48/XI65/XI5/MM1 N_XI48/XI65/NET21_XI48/XI65/XI5/MM1_d
+ N_XI48/XI65/NET52_XI48/XI65/XI5/MM1_g N_VSS_XI48/XI65/XI5/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI48/XI65/XI6/MM1 N_XI48/XI65/NET48_XI48/XI65/XI6/MM1_d
+ N_XI48/XI65/NET21_XI48/XI65/XI6/MM1_g N_VSS_XI48/XI65/XI6/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI48/XI64/XI5/MM1 N_XI48/XI64/NET21_XI48/XI64/XI5/MM1_d
+ N_XI48/XI64/NET52_XI48/XI64/XI5/MM1_g N_VSS_XI48/XI64/XI5/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI48/XI64/XI6/MM1 N_XI48/XI64/NET48_XI48/XI64/XI6/MM1_d
+ N_XI48/XI64/NET21_XI48/XI64/XI6/MM1_g N_VSS_XI48/XI64/XI6/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI48/XI60/XI6/MM1 N_XI48/XI60/NET48_XI48/XI60/XI6/MM1_d
+ N_XI48/XI60/NET21_XI48/XI60/XI6/MM1_g N_VSS_XI48/XI60/XI6/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI48/XI60/XI5/MM1 N_XI48/XI60/NET21_XI48/XI60/XI5/MM1_d
+ N_XI48/XI60/NET52_XI48/XI60/XI5/MM1_g N_VSS_XI48/XI60/XI5/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI48/XI61/XI5/MM1 N_XI48/XI61/NET21_XI48/XI61/XI5/MM1_d
+ N_XI48/XI61/NET52_XI48/XI61/XI5/MM1_g N_VSS_XI48/XI61/XI5/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI48/XI61/XI6/MM1 N_XI48/XI61/NET48_XI48/XI61/XI6/MM1_d
+ N_XI48/XI61/NET21_XI48/XI61/XI6/MM1_g N_VSS_XI48/XI61/XI6/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI48/XI62/XI6/MM1 N_XI48/XI62/NET48_XI48/XI62/XI6/MM1_d
+ N_XI48/XI62/NET21_XI48/XI62/XI6/MM1_g N_VSS_XI48/XI62/XI6/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI48/XI62/XI5/MM1 N_XI48/XI62/NET21_XI48/XI62/XI5/MM1_d
+ N_XI48/XI62/NET52_XI48/XI62/XI5/MM1_g N_VSS_XI48/XI62/XI5/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI48/XI63/XI5/MM1 N_XI48/XI63/NET21_XI48/XI63/XI5/MM1_d
+ N_XI48/XI63/NET52_XI48/XI63/XI5/MM1_g N_VSS_XI48/XI63/XI5/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI48/XI63/XI6/MM1 N_XI48/XI63/NET48_XI48/XI63/XI6/MM1_d
+ N_XI48/XI63/NET21_XI48/XI63/XI6/MM1_g N_VSS_XI48/XI63/XI6/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI32/XI9/XI13/MM1 N_XI32/XI9/NET21_XI32/XI9/XI13/MM1_d
+ N_XI32/XI9/NET52_XI32/XI9/XI13/MM1_g N_VSS_XI32/XI9/XI13/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI32/XI9/XI10/MM1 N_XI32/XI9/NET48_XI32/XI9/XI10/MM1_d
+ N_XI32/XI9/NET21_XI32/XI9/XI10/MM1_g N_VSS_XI32/XI9/XI10/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI32/XI8/XI13/MM1 N_XI32/XI8/NET21_XI32/XI8/XI13/MM1_d
+ N_XI32/XI8/NET52_XI32/XI8/XI13/MM1_g N_VSS_XI32/XI8/XI13/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI32/XI8/XI10/MM1 N_XI32/XI8/NET48_XI32/XI8/XI10/MM1_d
+ N_XI32/XI8/NET21_XI32/XI8/XI10/MM1_g N_VSS_XI32/XI8/XI10/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI32/XI7/XI13/MM1 N_XI32/XI7/NET21_XI32/XI7/XI13/MM1_d
+ N_XI32/XI7/NET52_XI32/XI7/XI13/MM1_g N_VSS_XI32/XI7/XI13/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI32/XI7/XI10/MM1 N_XI32/XI7/NET48_XI32/XI7/XI10/MM1_d
+ N_XI32/XI7/NET21_XI32/XI7/XI10/MM1_g N_VSS_XI32/XI7/XI10/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI42/XI519/XI72/XI20/MM5 N_XI42/XI519/NET113_XI42/XI519/XI72/XI20/MM5_d
+ N_NET128_XI42/XI519/XI72/XI20/MM5_g N_VSS_XI42/XI519/XI72/XI20/MM5_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13
+ AS=2.397e-13 PD=7.2e-07 PS=1.49e-06
mXI42/XI519/XI73/XI20/MM5 N_XI42/XI519/NET31_XI42/XI519/XI73/XI20/MM5_d
+ N_NET142_XI42/XI519/XI73/XI20/MM5_g N_VSS_XI42/XI519/XI73/XI20/MM5_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13
+ AS=2.397e-13 PD=7.2e-07 PS=1.49e-06
mXI48/XI74/XI3/MM1 N_NET136_XI48/XI74/XI3/MM1_d N_NET135_XI48/XI74/XI3/MM1_g
+ N_VSS_XI48/XI74/XI3/MM1_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=5e-07 AD=2.55e-13 AS=2.85e-13 PD=1.52e-06 PS=1.64e-06
mXI48/XI73/XI3/MM1 N_NET138_XI48/XI73/XI3/MM1_d N_NET137_XI48/XI73/XI3/MM1_g
+ N_VSS_XI48/XI73/XI3/MM1_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=5e-07 AD=2.55e-13 AS=2.85e-13 PD=1.52e-06 PS=1.64e-06
mXI48/XI72/XI3/MM1 N_NET140_XI48/XI72/XI3/MM1_d N_NET139_XI48/XI72/XI3/MM1_g
+ N_VSS_XI48/XI72/XI3/MM1_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=5e-07 AD=2.55e-13 AS=2.85e-13 PD=1.52e-06 PS=1.64e-06
mXI42/XI519/XI72/XI20/MM4 N_XI42/XI519/NET113_XI42/XI519/XI72/XI20/MM4_d
+ N_NET129_XI42/XI519/XI72/XI20/MM4_g N_VSS_XI42/XI519/XI72/XI20/MM4_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13
+ AS=2.397e-13 PD=7.2e-07 PS=1.49e-06
mXI42/XI519/XI73/XI20/MM4 N_XI42/XI519/NET31_XI42/XI519/XI73/XI20/MM4_d
+ N_NET143_XI42/XI519/XI73/XI20/MM4_g N_VSS_XI42/XI519/XI73/XI20/MM4_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13
+ AS=2.397e-13 PD=7.2e-07 PS=1.49e-06
mXI56/MM1 N_NET90_XI56/MM1_d N_CLK_XI56/MM1_g N_VSS_XI56/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI58/XI164/XI0/MM1 N_XI58/XI164/NET10_XI58/XI164/XI0/MM1_d
+ N_CLK_XI58/XI164/XI0/MM1_g N_VSS_XI58/XI164/XI0/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
mXI58/XI164/XI0/MM1@2 N_XI58/XI164/NET10_XI58/XI164/XI0/MM1@2_d
+ N_CLK_XI58/XI164/XI0/MM1@2_g N_VSS_XI58/XI164/XI0/MM1@2_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
mXI58/XI164/XI1/MM1 N_NET069_XI58/XI164/XI1/MM1_d
+ N_XI58/XI164/NET10_XI58/XI164/XI1/MM1_g N_VSS_XI58/XI164/XI1/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
mXI58/XI164/XI1/MM1@2 N_NET069_XI58/XI164/XI1/MM1@2_d
+ N_XI58/XI164/NET10_XI58/XI164/XI1/MM1@2_g N_VSS_XI58/XI164/XI1/MM1@2_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
mXI58/XI162/XI0/MM1 N_XI58/XI162/NET8_XI58/XI162/XI0/MM1_d
+ N_NET069_XI58/XI162/XI0/MM1_g N_VSS_XI58/XI162/XI0/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI58/XI162/XI1/MM1 N_XI58/NET086_XI58/XI162/XI1/MM1_d
+ N_XI58/XI162/NET8_XI58/XI162/XI1/MM1_g N_VSS_XI58/XI162/XI1/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI58/XI86/XI0/MM1 N_XI58/XI86/NET8_XI58/XI86/XI0/MM1_d
+ N_XI58/NET086_XI58/XI86/XI0/MM1_g N_VSS_XI58/XI86/XI0/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI58/XI86/XI1/MM1 N_XI58/NET30_XI58/XI86/XI1/MM1_d
+ N_XI58/XI86/NET8_XI58/XI86/XI1/MM1_g N_VSS_XI58/XI86/XI1/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI58/XI99/XI0/MM1 N_XI58/XI99/NET8_XI58/XI99/XI0/MM1_d
+ N_XI58/NET30_XI58/XI99/XI0/MM1_g N_VSS_XI58/XI99/XI0/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI58/XI99/XI1/MM1 N_XI58/NET039_XI58/XI99/XI1/MM1_d
+ N_XI58/XI99/NET8_XI58/XI99/XI1/MM1_g N_VSS_XI58/XI99/XI1/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI58/XI149/XI0/MM1 N_XI58/XI149/NET8_XI58/XI149/XI0/MM1_d
+ N_XI58/NET039_XI58/XI149/XI0/MM1_g N_VSS_XI58/XI149/XI0/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI58/XI149/XI1/MM1 N_XI58/NET081_XI58/XI149/XI1/MM1_d
+ N_XI58/XI149/NET8_XI58/XI149/XI1/MM1_g N_VSS_XI58/XI149/XI1/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI58/XI101/XI0/MM1 N_XI58/XI101/NET8_XI58/XI101/XI0/MM1_d
+ N_XI58/NET081_XI58/XI101/XI0/MM1_g N_VSS_XI58/XI101/XI0/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI58/XI101/XI1/MM1 N_NET070_XI58/XI101/XI1/MM1_d
+ N_XI58/XI101/NET8_XI58/XI101/XI1/MM1_g N_VSS_XI58/XI101/XI1/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI58/XI179/XI0/MM1 N_XI58/XI179/NET10_XI58/XI179/XI0/MM1_d
+ N_NET070_XI58/XI179/XI0/MM1_g N_VSS_XI58/XI179/XI0/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.65e-06 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI58/XI179/XI1/MM1 N_XI58/NET068_XI58/XI179/XI1/MM1_d
+ N_XI58/XI179/NET10_XI58/XI179/XI1/MM1_g N_VSS_XI58/XI179/XI1/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.65e-06 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI58/XI181/XI0/MM1 N_XI58/XI181/NET10_XI58/XI181/XI0/MM1_d
+ N_XI58/NET068_XI58/XI181/XI0/MM1_g N_VSS_XI58/XI181/XI0/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.65e-06 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI58/XI181/XI1/MM1 N_XI58/NET033_XI58/XI181/XI1/MM1_d
+ N_XI58/XI181/NET10_XI58/XI181/XI1/MM1_g N_VSS_XI58/XI181/XI1/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.65e-06 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI58/XI182/XI0/MM1 N_XI58/XI182/NET8_XI58/XI182/XI0/MM1_d
+ N_XI58/NET033_XI58/XI182/XI0/MM1_g N_VSS_XI58/XI182/XI0/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI58/XI182/XI1/MM1 N_XI58/NET049_XI58/XI182/XI1/MM1_d
+ N_XI58/XI182/NET8_XI58/XI182/XI1/MM1_g N_VSS_XI58/XI182/XI1/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI58/XI183/XI0/MM1 N_XI58/XI183/NET8_XI58/XI183/XI0/MM1_d
+ N_XI58/NET049_XI58/XI183/XI0/MM1_g N_VSS_XI58/XI183/XI0/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI58/XI183/XI1/MM1 N_NET068_XI58/XI183/XI1/MM1_d
+ N_XI58/XI183/NET8_XI58/XI183/XI1/MM1_g N_VSS_XI58/XI183/XI1/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI48/XI66/MM6 N_XI48/XI66/NET44_XI48/XI66/MM6_d N_CLK_XI48/XI66/MM6_g
+ N_XI48/XI66/NET21_XI48/XI66/MM6_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI48/XI66/MM7 N_XI48/XI66/NET059_XI48/XI66/MM7_d N_NET90_XI48/XI66/MM7_g
+ N_XI48/XI66/NET44_XI48/XI66/MM7_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI48/XI65/MM6 N_XI48/XI65/NET44_XI48/XI65/MM6_d N_CLK_XI48/XI65/MM6_g
+ N_XI48/XI65/NET21_XI48/XI65/MM6_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI48/XI65/MM7 N_XI48/XI65/NET059_XI48/XI65/MM7_d N_NET90_XI48/XI65/MM7_g
+ N_XI48/XI65/NET44_XI48/XI65/MM7_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI48/XI64/MM6 N_XI48/XI64/NET44_XI48/XI64/MM6_d N_CLK_XI48/XI64/MM6_g
+ N_XI48/XI64/NET21_XI48/XI64/MM6_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI48/XI64/MM7 N_XI48/XI64/NET059_XI48/XI64/MM7_d N_NET90_XI48/XI64/MM7_g
+ N_XI48/XI64/NET44_XI48/XI64/MM7_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI48/XI60/MM7 N_XI48/XI60/NET059_XI48/XI60/MM7_d N_NET90_XI48/XI60/MM7_g
+ N_XI48/XI60/NET44_XI48/XI60/MM7_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI48/XI60/MM6 N_XI48/XI60/NET44_XI48/XI60/MM6_d N_CLK_XI48/XI60/MM6_g
+ N_XI48/XI60/NET21_XI48/XI60/MM6_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI48/XI61/MM6 N_XI48/XI61/NET44_XI48/XI61/MM6_d N_CLK_XI48/XI61/MM6_g
+ N_XI48/XI61/NET21_XI48/XI61/MM6_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI48/XI61/MM7 N_XI48/XI61/NET059_XI48/XI61/MM7_d N_NET90_XI48/XI61/MM7_g
+ N_XI48/XI61/NET44_XI48/XI61/MM7_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI48/XI62/MM7 N_XI48/XI62/NET059_XI48/XI62/MM7_d N_NET90_XI48/XI62/MM7_g
+ N_XI48/XI62/NET44_XI48/XI62/MM7_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI48/XI62/MM6 N_XI48/XI62/NET44_XI48/XI62/MM6_d N_CLK_XI48/XI62/MM6_g
+ N_XI48/XI62/NET21_XI48/XI62/MM6_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI48/XI63/MM6 N_XI48/XI63/NET44_XI48/XI63/MM6_d N_CLK_XI48/XI63/MM6_g
+ N_XI48/XI63/NET21_XI48/XI63/MM6_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI48/XI63/MM7 N_XI48/XI63/NET059_XI48/XI63/MM7_d N_NET90_XI48/XI63/MM7_g
+ N_XI48/XI63/NET44_XI48/XI63/MM7_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI32/XI9/MM6 N_XI32/XI9/NET44_XI32/XI9/MM6_d N_CLK_XI32/XI9/MM6_g
+ N_XI32/XI9/NET21_XI32/XI9/MM6_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI32/XI9/MM7 N_NET434_XI32/XI9/MM7_d N_NET90_XI32/XI9/MM7_g
+ N_XI32/XI9/NET44_XI32/XI9/MM7_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI32/XI8/MM6 N_XI32/XI8/NET44_XI32/XI8/MM6_d N_CLK_XI32/XI8/MM6_g
+ N_XI32/XI8/NET21_XI32/XI8/MM6_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI32/XI8/MM7 N_NET435_XI32/XI8/MM7_d N_NET90_XI32/XI8/MM7_g
+ N_XI32/XI8/NET44_XI32/XI8/MM7_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI32/XI7/MM6 N_XI32/XI7/NET44_XI32/XI7/MM6_d N_CLK_XI32/XI7/MM6_g
+ N_XI32/XI7/NET21_XI32/XI7/MM6_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI32/XI7/MM7 N_NET436_XI32/XI7/MM7_d N_NET90_XI32/XI7/MM7_g
+ N_XI32/XI7/NET44_XI32/XI7/MM7_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI42/XI519/XI72/XI19/MM5 N_XI42/XI519/NET112_XI42/XI519/XI72/XI19/MM5_d
+ N_NET127_XI42/XI519/XI72/XI19/MM5_g N_VSS_XI42/XI519/XI72/XI19/MM5_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13
+ AS=2.397e-13 PD=7.2e-07 PS=1.49e-06
mXI42/XI519/XI73/XI19/MM5 N_XI42/XI519/NET104_XI42/XI519/XI73/XI19/MM5_d
+ N_NET141_XI42/XI519/XI73/XI19/MM5_g N_VSS_XI42/XI519/XI73/XI19/MM5_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13
+ AS=2.397e-13 PD=7.2e-07 PS=1.49e-06
mXI48/XI66/XI7/MM1 N_XI48/NET0110_XI48/XI66/XI7/MM1_d
+ N_XI48/XI66/NET44_XI48/XI66/XI7/MM1_g N_VSS_XI48/XI66/XI7/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI48/XI66/XI8/MM1 N_XI48/XI66/NET059_XI48/XI66/XI8/MM1_d
+ N_XI48/NET0110_XI48/XI66/XI8/MM1_g N_VSS_XI48/XI66/XI8/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI48/XI65/XI7/MM1 N_XI48/NET098_XI48/XI65/XI7/MM1_d
+ N_XI48/XI65/NET44_XI48/XI65/XI7/MM1_g N_VSS_XI48/XI65/XI7/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI48/XI65/XI8/MM1 N_XI48/XI65/NET059_XI48/XI65/XI8/MM1_d
+ N_XI48/NET098_XI48/XI65/XI8/MM1_g N_VSS_XI48/XI65/XI8/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI48/XI64/XI7/MM1 N_XI48/NET0116_XI48/XI64/XI7/MM1_d
+ N_XI48/XI64/NET44_XI48/XI64/XI7/MM1_g N_VSS_XI48/XI64/XI7/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI48/XI64/XI8/MM1 N_XI48/XI64/NET059_XI48/XI64/XI8/MM1_d
+ N_XI48/NET0116_XI48/XI64/XI8/MM1_g N_VSS_XI48/XI64/XI8/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI48/XI60/XI8/MM1 N_XI48/XI60/NET059_XI48/XI60/XI8/MM1_d
+ N_XI48/NET0122_XI48/XI60/XI8/MM1_g N_VSS_XI48/XI60/XI8/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI48/XI60/XI7/MM1 N_XI48/NET0122_XI48/XI60/XI7/MM1_d
+ N_XI48/XI60/NET44_XI48/XI60/XI7/MM1_g N_VSS_XI48/XI60/XI7/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI48/XI61/XI7/MM1 N_XI48/NET0134_XI48/XI61/XI7/MM1_d
+ N_XI48/XI61/NET44_XI48/XI61/XI7/MM1_g N_VSS_XI48/XI61/XI7/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI48/XI61/XI8/MM1 N_XI48/XI61/NET059_XI48/XI61/XI8/MM1_d
+ N_XI48/NET0134_XI48/XI61/XI8/MM1_g N_VSS_XI48/XI61/XI8/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI48/XI62/XI8/MM1 N_XI48/XI62/NET059_XI48/XI62/XI8/MM1_d
+ N_XI48/NET0128_XI48/XI62/XI8/MM1_g N_VSS_XI48/XI62/XI8/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI48/XI62/XI7/MM1 N_XI48/NET0128_XI48/XI62/XI7/MM1_d
+ N_XI48/XI62/NET44_XI48/XI62/XI7/MM1_g N_VSS_XI48/XI62/XI7/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI48/XI63/XI7/MM1 N_XI48/NET0104_XI48/XI63/XI7/MM1_d
+ N_XI48/XI63/NET44_XI48/XI63/XI7/MM1_g N_VSS_XI48/XI63/XI7/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI48/XI63/XI8/MM1 N_XI48/XI63/NET059_XI48/XI63/XI8/MM1_d
+ N_XI48/NET0104_XI48/XI63/XI8/MM1_g N_VSS_XI48/XI63/XI8/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI32/XI9/XI12/MM1 N_NET437_XI32/XI9/XI12/MM1_d
+ N_XI32/XI9/NET44_XI32/XI9/XI12/MM1_g N_VSS_XI32/XI9/XI12/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI32/XI9/XI11/MM1 N_NET434_XI32/XI9/XI11/MM1_d N_NET437_XI32/XI9/XI11/MM1_g
+ N_VSS_XI32/XI9/XI11/MM1_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI32/XI8/XI12/MM1 N_NET438_XI32/XI8/XI12/MM1_d
+ N_XI32/XI8/NET44_XI32/XI8/XI12/MM1_g N_VSS_XI32/XI8/XI12/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI32/XI8/XI11/MM1 N_NET435_XI32/XI8/XI11/MM1_d N_NET438_XI32/XI8/XI11/MM1_g
+ N_VSS_XI32/XI8/XI11/MM1_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI32/XI7/XI12/MM1 N_NET439_XI32/XI7/XI12/MM1_d
+ N_XI32/XI7/NET44_XI32/XI7/XI12/MM1_g N_VSS_XI32/XI7/XI12/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI32/XI7/XI11/MM1 N_NET436_XI32/XI7/XI11/MM1_d N_NET439_XI32/XI7/XI11/MM1_g
+ N_VSS_XI32/XI7/XI11/MM1_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI42/XI519/XI72/XI19/MM4 N_XI42/XI519/NET112_XI42/XI519/XI72/XI19/MM4_d
+ N_NET130_XI42/XI519/XI72/XI19/MM4_g N_VSS_XI42/XI519/XI72/XI19/MM4_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13
+ AS=2.397e-13 PD=7.2e-07 PS=1.49e-06
mXI42/XI519/XI73/XI19/MM4 N_XI42/XI519/NET104_XI42/XI519/XI73/XI19/MM4_d
+ N_NET126_XI42/XI519/XI73/XI19/MM4_g N_VSS_XI42/XI519/XI73/XI19/MM4_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13
+ AS=2.397e-13 PD=7.2e-07 PS=1.49e-06
mXI30/XI67/MM5 N_XI30/XI67/NET7_XI30/XI67/MM5_d N_NET437_XI30/XI67/MM5_g
+ N_VSS_XI30/XI67/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI30/XI67/MM4 N_XI30/XI67/NET11_XI30/XI67/MM4_d N_NET438_XI30/XI67/MM4_g
+ N_XI30/XI67/NET7_XI30/XI67/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18
+ L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI30/XI67/MM3 N_NET470_XI30/XI67/MM3_d N_NET439_XI30/XI67/MM3_g
+ N_XI30/XI67/NET11_XI30/XI67/MM3_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18
+ L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI30/XI69/MM5 N_XI30/XI69/NET7_XI30/XI69/MM5_d N_NET437_XI30/XI69/MM5_g
+ N_VSS_XI30/XI69/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI30/XI69/MM4 N_XI30/XI69/NET11_XI30/XI69/MM4_d N_NET435_XI30/XI69/MM4_g
+ N_XI30/XI69/NET7_XI30/XI69/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18
+ L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI30/XI69/MM3 N_NET468_XI30/XI69/MM3_d N_NET439_XI30/XI69/MM3_g
+ N_XI30/XI69/NET11_XI30/XI69/MM3_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18
+ L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI30/XI71/MM5 N_XI30/XI71/NET7_XI30/XI71/MM5_d N_NET437_XI30/XI71/MM5_g
+ N_VSS_XI30/XI71/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI30/XI71/MM4 N_XI30/XI71/NET11_XI30/XI71/MM4_d N_NET438_XI30/XI71/MM4_g
+ N_XI30/XI71/NET7_XI30/XI71/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18
+ L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI30/XI71/MM3 N_NET466_XI30/XI71/MM3_d N_NET436_XI30/XI71/MM3_g
+ N_XI30/XI71/NET11_XI30/XI71/MM3_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18
+ L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI30/XI73/MM5 N_XI30/XI73/NET7_XI30/XI73/MM5_d N_NET437_XI30/XI73/MM5_g
+ N_VSS_XI30/XI73/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI30/XI73/MM4 N_XI30/XI73/NET11_XI30/XI73/MM4_d N_NET435_XI30/XI73/MM4_g
+ N_XI30/XI73/NET7_XI30/XI73/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18
+ L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI30/XI73/MM3 N_NET464_XI30/XI73/MM3_d N_NET436_XI30/XI73/MM3_g
+ N_XI30/XI73/NET11_XI30/XI73/MM3_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18
+ L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI30/XI68/MM5 N_XI30/XI68/NET7_XI30/XI68/MM5_d N_NET434_XI30/XI68/MM5_g
+ N_VSS_XI30/XI68/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI30/XI68/MM4 N_XI30/XI68/NET11_XI30/XI68/MM4_d N_NET438_XI30/XI68/MM4_g
+ N_XI30/XI68/NET7_XI30/XI68/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18
+ L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI30/XI68/MM3 N_NET469_XI30/XI68/MM3_d N_NET439_XI30/XI68/MM3_g
+ N_XI30/XI68/NET11_XI30/XI68/MM3_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18
+ L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI30/XI70/MM5 N_XI30/XI70/NET7_XI30/XI70/MM5_d N_NET434_XI30/XI70/MM5_g
+ N_VSS_XI30/XI70/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI30/XI70/MM4 N_XI30/XI70/NET11_XI30/XI70/MM4_d N_NET435_XI30/XI70/MM4_g
+ N_XI30/XI70/NET7_XI30/XI70/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18
+ L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI30/XI70/MM3 N_NET467_XI30/XI70/MM3_d N_NET439_XI30/XI70/MM3_g
+ N_XI30/XI70/NET11_XI30/XI70/MM3_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18
+ L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI30/XI72/MM5 N_XI30/XI72/NET7_XI30/XI72/MM5_d N_NET434_XI30/XI72/MM5_g
+ N_VSS_XI30/XI72/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI30/XI72/MM4 N_XI30/XI72/NET11_XI30/XI72/MM4_d N_NET438_XI30/XI72/MM4_g
+ N_XI30/XI72/NET7_XI30/XI72/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18
+ L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI30/XI72/MM3 N_NET465_XI30/XI72/MM3_d N_NET436_XI30/XI72/MM3_g
+ N_XI30/XI72/NET11_XI30/XI72/MM3_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18
+ L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI30/XI74/MM5 N_XI30/XI74/NET7_XI30/XI74/MM5_d N_NET434_XI30/XI74/MM5_g
+ N_VSS_XI30/XI74/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI30/XI74/MM4 N_XI30/XI74/NET11_XI30/XI74/MM4_d N_NET435_XI30/XI74/MM4_g
+ N_XI30/XI74/NET7_XI30/XI74/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18
+ L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI30/XI74/MM3 N_NET463_XI30/XI74/MM3_d N_NET436_XI30/XI74/MM3_g
+ N_XI30/XI74/NET11_XI30/XI74/MM3_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18
+ L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI42/XI652/XI0/MM1 N_XI42/XI652/NET8_XI42/XI652/XI0/MM1_d
+ N_XI42/NET01023_XI42/XI652/XI0/MM1_g N_VSS_XI42/XI652/XI0/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI48/XI74/XI2/MM3 N_XI48/XI74/XI2/NET13_XI48/XI74/XI2/MM3_d
+ N_XI48/NET0110_XI48/XI74/XI2/MM3_g N_VSS_XI48/XI74/XI2/MM3_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13
+ AS=2.397e-13 PD=7.2e-07 PS=1.49e-06
mXI48/XI73/XI2/MM3 N_XI48/XI73/XI2/NET13_XI48/XI73/XI2/MM3_d
+ N_XI48/NET098_XI48/XI73/XI2/MM3_g N_VSS_XI48/XI73/XI2/MM3_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13
+ AS=2.397e-13 PD=7.2e-07 PS=1.49e-06
mXI48/XI72/XI2/MM3 N_XI48/XI72/XI2/NET13_XI48/XI72/XI2/MM3_d
+ N_XI48/NET0116_XI48/XI72/XI2/MM3_g N_VSS_XI48/XI72/XI2/MM3_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13
+ AS=2.397e-13 PD=7.2e-07 PS=1.49e-06
mXI42/XI519/XI72/XI18/MM5 N_XI42/XI519/NET111_XI42/XI519/XI72/XI18/MM5_d
+ N_NET128_XI42/XI519/XI72/XI18/MM5_g N_VSS_XI42/XI519/XI72/XI18/MM5_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13
+ AS=2.397e-13 PD=7.2e-07 PS=1.49e-06
mXI42/XI519/XI73/XI18/MM5 N_XI42/XI519/NET103_XI42/XI519/XI73/XI18/MM5_d
+ N_NET142_XI42/XI519/XI73/XI18/MM5_g N_VSS_XI42/XI519/XI73/XI18/MM5_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13
+ AS=2.397e-13 PD=7.2e-07 PS=1.49e-06
mXI48/XI74/XI2/MM2 N_NET135_XI48/XI74/XI2/MM2_d N_NET069_XI48/XI74/XI2/MM2_g
+ N_XI48/XI74/XI2/NET13_XI48/XI74/XI2/MM2_s N_VSS_XI42/XI519/XI72/XI21/MM5_b
+ N_18 L=1.8e-07 W=4.7e-07 AD=2.397e-13 AS=1.692e-13 PD=1.49e-06 PS=7.2e-07
mXI48/XI73/XI2/MM2 N_NET137_XI48/XI73/XI2/MM2_d N_NET069_XI48/XI73/XI2/MM2_g
+ N_XI48/XI73/XI2/NET13_XI48/XI73/XI2/MM2_s N_VSS_XI42/XI519/XI72/XI21/MM5_b
+ N_18 L=1.8e-07 W=4.7e-07 AD=2.397e-13 AS=1.692e-13 PD=1.49e-06 PS=7.2e-07
mXI48/XI72/XI2/MM2 N_NET139_XI48/XI72/XI2/MM2_d N_NET069_XI48/XI72/XI2/MM2_g
+ N_XI48/XI72/XI2/NET13_XI48/XI72/XI2/MM2_s N_VSS_XI42/XI519/XI72/XI21/MM5_b
+ N_18 L=1.8e-07 W=4.7e-07 AD=2.397e-13 AS=1.692e-13 PD=1.49e-06 PS=7.2e-07
mXI42/XI519/XI72/XI18/MM4 N_XI42/XI519/NET111_XI42/XI519/XI72/XI18/MM4_d
+ N_NET130_XI42/XI519/XI72/XI18/MM4_g N_VSS_XI42/XI519/XI72/XI18/MM4_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13
+ AS=2.397e-13 PD=7.2e-07 PS=1.49e-06
mXI42/XI519/XI73/XI18/MM4 N_XI42/XI519/NET103_XI42/XI519/XI73/XI18/MM4_d
+ N_NET126_XI42/XI519/XI73/XI18/MM4_g N_VSS_XI42/XI519/XI73/XI18/MM4_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13
+ AS=2.397e-13 PD=7.2e-07 PS=1.49e-06
mXI42/XI652/XI1/MM1 N_NET0133_XI42/XI652/XI1/MM1_d
+ N_XI42/XI652/NET8_XI42/XI652/XI1/MM1_g N_VSS_XI42/XI652/XI1/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI48/XI68/XI2/MM3 N_XI48/XI68/XI2/NET13_XI48/XI68/XI2/MM3_d
+ N_XI48/NET0122_XI48/XI68/XI2/MM3_g N_VSS_XI48/XI68/XI2/MM3_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13
+ AS=2.397e-13 PD=7.2e-07 PS=1.49e-06
mXI48/XI68/XI2/MM2 N_NET129_XI48/XI68/XI2/MM2_d N_NET069_XI48/XI68/XI2/MM2_g
+ N_XI48/XI68/XI2/NET13_XI48/XI68/XI2/MM2_s N_VSS_XI42/XI519/XI72/XI21/MM5_b
+ N_18 L=1.8e-07 W=4.7e-07 AD=2.397e-13 AS=1.692e-13 PD=1.49e-06 PS=7.2e-07
mXI48/XI70/XI2/MM3 N_XI48/XI70/XI2/NET13_XI48/XI70/XI2/MM3_d
+ N_XI48/NET0128_XI48/XI70/XI2/MM3_g N_VSS_XI48/XI70/XI2/MM3_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13
+ AS=2.397e-13 PD=7.2e-07 PS=1.49e-06
mXI48/XI70/XI2/MM2 N_NET143_XI48/XI70/XI2/MM2_d N_NET069_XI48/XI70/XI2/MM2_g
+ N_XI48/XI70/XI2/NET13_XI48/XI70/XI2/MM2_s N_VSS_XI42/XI519/XI72/XI21/MM5_b
+ N_18 L=1.8e-07 W=4.7e-07 AD=2.397e-13 AS=1.692e-13 PD=1.49e-06 PS=7.2e-07
mXI48/XI69/XI2/MM2 N_NET127_XI48/XI69/XI2/MM2_d N_NET069_XI48/XI69/XI2/MM2_g
+ N_XI48/XI69/XI2/NET13_XI48/XI69/XI2/MM2_s N_VSS_XI42/XI519/XI72/XI21/MM5_b
+ N_18 L=1.8e-07 W=4.7e-07 AD=2.397e-13 AS=1.692e-13 PD=1.49e-06 PS=7.2e-07
mXI48/XI69/XI2/MM3 N_XI48/XI69/XI2/NET13_XI48/XI69/XI2/MM3_d
+ N_XI48/NET0134_XI48/XI69/XI2/MM3_g N_VSS_XI48/XI69/XI2/MM3_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13
+ AS=2.397e-13 PD=7.2e-07 PS=1.49e-06
mXI48/XI71/XI2/MM2 N_NET141_XI48/XI71/XI2/MM2_d N_NET069_XI48/XI71/XI2/MM2_g
+ N_XI48/XI71/XI2/NET13_XI48/XI71/XI2/MM2_s N_VSS_XI42/XI519/XI72/XI21/MM5_b
+ N_18 L=1.8e-07 W=4.7e-07 AD=2.397e-13 AS=1.692e-13 PD=1.49e-06 PS=7.2e-07
mXI48/XI71/XI2/MM3 N_XI48/XI71/XI2/NET13_XI48/XI71/XI2/MM3_d
+ N_XI48/NET0104_XI48/XI71/XI2/MM3_g N_VSS_XI48/XI71/XI2/MM3_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13
+ AS=2.397e-13 PD=7.2e-07 PS=1.49e-06
mXI48/XI68/XI3/MM1 N_NET130_XI48/XI68/XI3/MM1_d N_NET129_XI48/XI68/XI3/MM1_g
+ N_VSS_XI48/XI68/XI3/MM1_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI48/XI69/XI3/MM1 N_NET128_XI48/XI69/XI3/MM1_d N_NET127_XI48/XI69/XI3/MM1_g
+ N_VSS_XI48/XI69/XI3/MM1_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI48/XI70/XI3/MM1 N_NET126_XI48/XI70/XI3/MM1_d N_NET143_XI48/XI70/XI3/MM1_g
+ N_VSS_XI48/XI70/XI3/MM1_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI48/XI71/XI3/MM1 N_NET142_XI48/XI71/XI3/MM1_d N_NET141_XI48/XI71/XI3/MM1_g
+ N_VSS_XI48/XI71/XI3/MM1_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI54/XI0/XI10/MM4 N_DOUT<0>_XI54/XI0/XI10/MM4_d
+ N_XI54/NET10_XI54/XI0/XI10/MM4_g N_VSS_XI54/XI0/XI10/MM4_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=1.68025e-13
+ AS=2.3265e-13 PD=7.15e-07 PS=1.46e-06
mXI54/XI0/XI9/MM4 N_XI54/NET10_XI54/XI0/XI9/MM4_d
+ N_XI54/XI0/NET10_XI54/XI0/XI9/MM4_g N_VSS_XI54/XI0/XI9/MM4_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=1.68025e-13
+ AS=2.3265e-13 PD=7.15e-07 PS=1.46e-06
mXI54/XI0/XI10/MM5 N_DOUT<0>_XI54/XI0/XI10/MM5_d
+ N_XI54/XI0/NET9_XI54/XI0/XI10/MM5_g N_VSS_XI54/XI0/XI10/MM5_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=1.68025e-13
+ AS=2.303e-13 PD=7.15e-07 PS=1.45e-06
mXI54/XI0/XI9/MM5 N_XI54/NET10_XI54/XI0/XI9/MM5_d N_DOUT<0>_XI54/XI0/XI9/MM5_g
+ N_VSS_XI54/XI0/XI9/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.68025e-13 AS=2.303e-13 PD=7.15e-07 PS=1.45e-06
mXI54/XI0/XI8/XI2/MM1 N_XI54/XI0/NET9_XI54/XI0/XI8/XI2/MM1_d
+ N_XI54/XI0/XI8/NET12_XI54/XI0/XI8/XI2/MM1_g N_VSS_XI54/XI0/XI8/XI2/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13
+ AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI54/XI0/XI7/XI2/MM1 N_XI54/XI0/NET10_XI54/XI0/XI7/XI2/MM1_d
+ N_XI54/XI0/XI7/NET12_XI54/XI0/XI7/XI2/MM1_g N_VSS_XI54/XI0/XI7/XI2/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13
+ AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI42/XI519/XI86/MM2 N_XI42/NET780_XI42/XI519/XI86/MM2_d
+ N_XI42/XI519/NET114_XI42/XI519/XI86/MM2_g
+ N_XI42/XI519/XI86/NET13_XI42/XI519/XI86/MM2_s N_VSS_XI42/XI519/XI72/XI21/MM5_b
+ N_18 L=1.8e-07 W=4.7e-07 AD=2.397e-13 AS=1.692e-13 PD=1.49e-06 PS=7.2e-07
mXI42/XI519/XI86/MM3 N_XI42/XI519/XI86/NET13_XI42/XI519/XI86/MM3_d
+ N_XI42/XI519/NET36_XI42/XI519/XI86/MM3_g N_VSS_XI42/XI519/XI86/MM3_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13
+ AS=2.679e-13 PD=7.2e-07 PS=1.61e-06
mXI42/XI519/XI87/MM2 N_XI42/NET781_XI42/XI519/XI87/MM2_d
+ N_XI42/XI519/NET114_XI42/XI519/XI87/MM2_g
+ N_XI42/XI519/XI87/NET13_XI42/XI519/XI87/MM2_s N_VSS_XI42/XI519/XI72/XI21/MM5_b
+ N_18 L=1.8e-07 W=4.7e-07 AD=2.397e-13 AS=1.692e-13 PD=1.49e-06 PS=7.2e-07
mXI42/XI519/XI87/MM3 N_XI42/XI519/XI87/NET13_XI42/XI519/XI87/MM3_d
+ N_XI42/XI519/NET31_XI42/XI519/XI87/MM3_g N_VSS_XI42/XI519/XI87/MM3_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13
+ AS=2.679e-13 PD=7.2e-07 PS=1.61e-06
mXI42/XI519/XI88/MM2 N_XI42/NET782_XI42/XI519/XI88/MM2_d
+ N_XI42/XI519/NET114_XI42/XI519/XI88/MM2_g
+ N_XI42/XI519/XI88/NET13_XI42/XI519/XI88/MM2_s N_VSS_XI42/XI519/XI72/XI21/MM5_b
+ N_18 L=1.8e-07 W=4.7e-07 AD=2.397e-13 AS=1.692e-13 PD=1.49e-06 PS=7.2e-07
mXI42/XI519/XI88/MM3 N_XI42/XI519/XI88/NET13_XI42/XI519/XI88/MM3_d
+ N_XI42/XI519/NET104_XI42/XI519/XI88/MM3_g N_VSS_XI42/XI519/XI88/MM3_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13
+ AS=2.679e-13 PD=7.2e-07 PS=1.61e-06
mXI42/XI519/XI89/MM2 N_XI42/NET783_XI42/XI519/XI89/MM2_d
+ N_XI42/XI519/NET114_XI42/XI519/XI89/MM2_g
+ N_XI42/XI519/XI89/NET13_XI42/XI519/XI89/MM2_s N_VSS_XI42/XI519/XI72/XI21/MM5_b
+ N_18 L=1.8e-07 W=4.7e-07 AD=2.397e-13 AS=1.692e-13 PD=1.49e-06 PS=7.2e-07
mXI42/XI519/XI89/MM3 N_XI42/XI519/XI89/NET13_XI42/XI519/XI89/MM3_d
+ N_XI42/XI519/NET103_XI42/XI519/XI89/MM3_g N_VSS_XI42/XI519/XI89/MM3_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13
+ AS=2.679e-13 PD=7.2e-07 PS=1.61e-06
mXI42/XI519/XI82/MM2 N_XI42/NET784_XI42/XI519/XI82/MM2_d
+ N_XI42/XI519/NET113_XI42/XI519/XI82/MM2_g
+ N_XI42/XI519/XI82/NET13_XI42/XI519/XI82/MM2_s N_VSS_XI42/XI519/XI72/XI21/MM5_b
+ N_18 L=1.8e-07 W=4.7e-07 AD=2.397e-13 AS=1.692e-13 PD=1.49e-06 PS=7.2e-07
mXI42/XI519/XI82/MM3 N_XI42/XI519/XI82/NET13_XI42/XI519/XI82/MM3_d
+ N_XI42/XI519/NET36_XI42/XI519/XI82/MM3_g N_VSS_XI42/XI519/XI82/MM3_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13
+ AS=2.679e-13 PD=7.2e-07 PS=1.61e-06
mXI42/XI519/XI83/MM2 N_XI42/NET785_XI42/XI519/XI83/MM2_d
+ N_XI42/XI519/NET113_XI42/XI519/XI83/MM2_g
+ N_XI42/XI519/XI83/NET13_XI42/XI519/XI83/MM2_s N_VSS_XI42/XI519/XI72/XI21/MM5_b
+ N_18 L=1.8e-07 W=4.7e-07 AD=2.397e-13 AS=1.692e-13 PD=1.49e-06 PS=7.2e-07
mXI42/XI519/XI83/MM3 N_XI42/XI519/XI83/NET13_XI42/XI519/XI83/MM3_d
+ N_XI42/XI519/NET31_XI42/XI519/XI83/MM3_g N_VSS_XI42/XI519/XI83/MM3_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13
+ AS=2.679e-13 PD=7.2e-07 PS=1.61e-06
mXI42/XI519/XI84/MM2 N_XI42/NET786_XI42/XI519/XI84/MM2_d
+ N_XI42/XI519/NET113_XI42/XI519/XI84/MM2_g
+ N_XI42/XI519/XI84/NET13_XI42/XI519/XI84/MM2_s N_VSS_XI42/XI519/XI72/XI21/MM5_b
+ N_18 L=1.8e-07 W=4.7e-07 AD=2.397e-13 AS=1.692e-13 PD=1.49e-06 PS=7.2e-07
mXI42/XI519/XI84/MM3 N_XI42/XI519/XI84/NET13_XI42/XI519/XI84/MM3_d
+ N_XI42/XI519/NET104_XI42/XI519/XI84/MM3_g N_VSS_XI42/XI519/XI84/MM3_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13
+ AS=2.679e-13 PD=7.2e-07 PS=1.61e-06
mXI42/XI519/XI85/MM2 N_XI42/NET787_XI42/XI519/XI85/MM2_d
+ N_XI42/XI519/NET113_XI42/XI519/XI85/MM2_g
+ N_XI42/XI519/XI85/NET13_XI42/XI519/XI85/MM2_s N_VSS_XI42/XI519/XI72/XI21/MM5_b
+ N_18 L=1.8e-07 W=4.7e-07 AD=2.397e-13 AS=1.692e-13 PD=1.49e-06 PS=7.2e-07
mXI42/XI519/XI85/MM3 N_XI42/XI519/XI85/NET13_XI42/XI519/XI85/MM3_d
+ N_XI42/XI519/NET103_XI42/XI519/XI85/MM3_g N_VSS_XI42/XI519/XI85/MM3_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13
+ AS=2.679e-13 PD=7.2e-07 PS=1.61e-06
mXI42/XI519/XI78/MM2 N_XI42/NET788_XI42/XI519/XI78/MM2_d
+ N_XI42/XI519/NET112_XI42/XI519/XI78/MM2_g
+ N_XI42/XI519/XI78/NET13_XI42/XI519/XI78/MM2_s N_VSS_XI42/XI519/XI72/XI21/MM5_b
+ N_18 L=1.8e-07 W=4.7e-07 AD=2.397e-13 AS=1.692e-13 PD=1.49e-06 PS=7.2e-07
mXI42/XI519/XI78/MM3 N_XI42/XI519/XI78/NET13_XI42/XI519/XI78/MM3_d
+ N_XI42/XI519/NET36_XI42/XI519/XI78/MM3_g N_VSS_XI42/XI519/XI78/MM3_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13
+ AS=2.679e-13 PD=7.2e-07 PS=1.61e-06
mXI42/XI519/XI79/MM2 N_XI42/NET789_XI42/XI519/XI79/MM2_d
+ N_XI42/XI519/NET112_XI42/XI519/XI79/MM2_g
+ N_XI42/XI519/XI79/NET13_XI42/XI519/XI79/MM2_s N_VSS_XI42/XI519/XI72/XI21/MM5_b
+ N_18 L=1.8e-07 W=4.7e-07 AD=2.397e-13 AS=1.692e-13 PD=1.49e-06 PS=7.2e-07
mXI42/XI519/XI79/MM3 N_XI42/XI519/XI79/NET13_XI42/XI519/XI79/MM3_d
+ N_XI42/XI519/NET31_XI42/XI519/XI79/MM3_g N_VSS_XI42/XI519/XI79/MM3_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13
+ AS=2.679e-13 PD=7.2e-07 PS=1.61e-06
mXI42/XI519/XI80/MM2 N_XI42/NET790_XI42/XI519/XI80/MM2_d
+ N_XI42/XI519/NET112_XI42/XI519/XI80/MM2_g
+ N_XI42/XI519/XI80/NET13_XI42/XI519/XI80/MM2_s N_VSS_XI42/XI519/XI72/XI21/MM5_b
+ N_18 L=1.8e-07 W=4.7e-07 AD=2.397e-13 AS=1.692e-13 PD=1.49e-06 PS=7.2e-07
mXI42/XI519/XI80/MM3 N_XI42/XI519/XI80/NET13_XI42/XI519/XI80/MM3_d
+ N_XI42/XI519/NET104_XI42/XI519/XI80/MM3_g N_VSS_XI42/XI519/XI80/MM3_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13
+ AS=2.679e-13 PD=7.2e-07 PS=1.61e-06
mXI42/XI519/XI81/MM2 N_XI42/NET791_XI42/XI519/XI81/MM2_d
+ N_XI42/XI519/NET112_XI42/XI519/XI81/MM2_g
+ N_XI42/XI519/XI81/NET13_XI42/XI519/XI81/MM2_s N_VSS_XI42/XI519/XI72/XI21/MM5_b
+ N_18 L=1.8e-07 W=4.7e-07 AD=2.397e-13 AS=1.692e-13 PD=1.49e-06 PS=7.2e-07
mXI42/XI519/XI81/MM3 N_XI42/XI519/XI81/NET13_XI42/XI519/XI81/MM3_d
+ N_XI42/XI519/NET103_XI42/XI519/XI81/MM3_g N_VSS_XI42/XI519/XI81/MM3_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13
+ AS=2.679e-13 PD=7.2e-07 PS=1.61e-06
mXI42/XI519/XI74/MM2 N_XI42/NET792_XI42/XI519/XI74/MM2_d
+ N_XI42/XI519/NET111_XI42/XI519/XI74/MM2_g
+ N_XI42/XI519/XI74/NET13_XI42/XI519/XI74/MM2_s N_VSS_XI42/XI519/XI72/XI21/MM5_b
+ N_18 L=1.8e-07 W=4.7e-07 AD=2.397e-13 AS=1.692e-13 PD=1.49e-06 PS=7.2e-07
mXI42/XI519/XI74/MM3 N_XI42/XI519/XI74/NET13_XI42/XI519/XI74/MM3_d
+ N_XI42/XI519/NET36_XI42/XI519/XI74/MM3_g N_VSS_XI42/XI519/XI74/MM3_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13
+ AS=2.679e-13 PD=7.2e-07 PS=1.61e-06
mXI42/XI519/XI75/MM2 N_XI42/NET793_XI42/XI519/XI75/MM2_d
+ N_XI42/XI519/NET111_XI42/XI519/XI75/MM2_g
+ N_XI42/XI519/XI75/NET13_XI42/XI519/XI75/MM2_s N_VSS_XI42/XI519/XI72/XI21/MM5_b
+ N_18 L=1.8e-07 W=4.7e-07 AD=2.397e-13 AS=1.692e-13 PD=1.49e-06 PS=7.2e-07
mXI42/XI519/XI75/MM3 N_XI42/XI519/XI75/NET13_XI42/XI519/XI75/MM3_d
+ N_XI42/XI519/NET31_XI42/XI519/XI75/MM3_g N_VSS_XI42/XI519/XI75/MM3_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13
+ AS=2.679e-13 PD=7.2e-07 PS=1.61e-06
mXI42/XI519/XI76/MM2 N_XI42/NET794_XI42/XI519/XI76/MM2_d
+ N_XI42/XI519/NET111_XI42/XI519/XI76/MM2_g
+ N_XI42/XI519/XI76/NET13_XI42/XI519/XI76/MM2_s N_VSS_XI42/XI519/XI72/XI21/MM5_b
+ N_18 L=1.8e-07 W=4.7e-07 AD=2.397e-13 AS=1.692e-13 PD=1.49e-06 PS=7.2e-07
mXI42/XI519/XI76/MM3 N_XI42/XI519/XI76/NET13_XI42/XI519/XI76/MM3_d
+ N_XI42/XI519/NET104_XI42/XI519/XI76/MM3_g N_VSS_XI42/XI519/XI76/MM3_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13
+ AS=2.679e-13 PD=7.2e-07 PS=1.61e-06
mXI42/XI519/XI77/MM2 N_XI42/NET795_XI42/XI519/XI77/MM2_d
+ N_XI42/XI519/NET111_XI42/XI519/XI77/MM2_g
+ N_XI42/XI519/XI77/NET13_XI42/XI519/XI77/MM2_s N_VSS_XI42/XI519/XI72/XI21/MM5_b
+ N_18 L=1.8e-07 W=4.7e-07 AD=2.397e-13 AS=1.692e-13 PD=1.49e-06 PS=7.2e-07
mXI42/XI519/XI77/MM3 N_XI42/XI519/XI77/NET13_XI42/XI519/XI77/MM3_d
+ N_XI42/XI519/NET103_XI42/XI519/XI77/MM3_g N_VSS_XI42/XI519/XI77/MM3_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13
+ AS=2.679e-13 PD=7.2e-07 PS=1.61e-06
mXI42/XI520/XI12/MM16 N_XI42/NET801_XI42/XI520/XI12/MM16_d
+ N_NET140_XI42/XI520/XI12/MM16_g
+ N_XI42/XI520/XI12/NET034_XI42/XI520/XI12/MM16_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI42/XI520/XI12/MM17 N_XI42/XI520/XI12/NET034_XI42/XI520/XI12/MM17_d
+ N_NET138_XI42/XI520/XI12/MM17_g
+ N_XI42/XI520/XI12/NET048_XI42/XI520/XI12/MM17_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13
+ AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI42/XI520/XI12/MM18 N_XI42/XI520/XI12/NET048_XI42/XI520/XI12/MM18_d
+ N_NET136_XI42/XI520/XI12/MM18_g N_VSS_XI42/XI520/XI12/MM18_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13
+ AS=2.726e-13 PD=5.1e-07 PS=1.63e-06
mXI42/XI520/XI13/MM16 N_XI42/NET455_XI42/XI520/XI13/MM16_d
+ N_NET140_XI42/XI520/XI13/MM16_g
+ N_XI42/XI520/XI13/NET034_XI42/XI520/XI13/MM16_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI42/XI520/XI13/MM17 N_XI42/XI520/XI13/NET034_XI42/XI520/XI13/MM17_d
+ N_NET138_XI42/XI520/XI13/MM17_g
+ N_XI42/XI520/XI13/NET048_XI42/XI520/XI13/MM17_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13
+ AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI42/XI520/XI13/MM18 N_XI42/XI520/XI13/NET048_XI42/XI520/XI13/MM18_d
+ N_NET135_XI42/XI520/XI13/MM18_g N_VSS_XI42/XI520/XI13/MM18_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13
+ AS=2.726e-13 PD=5.1e-07 PS=1.63e-06
mXI42/XI520/XI14/MM16 N_XI42/NET803_XI42/XI520/XI14/MM16_d
+ N_NET140_XI42/XI520/XI14/MM16_g
+ N_XI42/XI520/XI14/NET034_XI42/XI520/XI14/MM16_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI42/XI520/XI14/MM17 N_XI42/XI520/XI14/NET034_XI42/XI520/XI14/MM17_d
+ N_NET137_XI42/XI520/XI14/MM17_g
+ N_XI42/XI520/XI14/NET048_XI42/XI520/XI14/MM17_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13
+ AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI42/XI520/XI14/MM18 N_XI42/XI520/XI14/NET048_XI42/XI520/XI14/MM18_d
+ N_NET136_XI42/XI520/XI14/MM18_g N_VSS_XI42/XI520/XI14/MM18_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13
+ AS=2.726e-13 PD=5.1e-07 PS=1.63e-06
mXI42/XI520/XI15/MM16 N_XI42/NET245_XI42/XI520/XI15/MM16_d
+ N_NET140_XI42/XI520/XI15/MM16_g
+ N_XI42/XI520/XI15/NET034_XI42/XI520/XI15/MM16_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI42/XI520/XI15/MM17 N_XI42/XI520/XI15/NET034_XI42/XI520/XI15/MM17_d
+ N_NET137_XI42/XI520/XI15/MM17_g
+ N_XI42/XI520/XI15/NET048_XI42/XI520/XI15/MM17_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13
+ AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI42/XI520/XI15/MM18 N_XI42/XI520/XI15/NET048_XI42/XI520/XI15/MM18_d
+ N_NET135_XI42/XI520/XI15/MM18_g N_VSS_XI42/XI520/XI15/MM18_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13
+ AS=2.726e-13 PD=5.1e-07 PS=1.63e-06
mXI42/XI520/XI16/MM16 N_XI42/NET802_XI42/XI520/XI16/MM16_d
+ N_NET139_XI42/XI520/XI16/MM16_g
+ N_XI42/XI520/XI16/NET034_XI42/XI520/XI16/MM16_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI42/XI520/XI16/MM17 N_XI42/XI520/XI16/NET034_XI42/XI520/XI16/MM17_d
+ N_NET138_XI42/XI520/XI16/MM17_g
+ N_XI42/XI520/XI16/NET048_XI42/XI520/XI16/MM17_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13
+ AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI42/XI520/XI16/MM18 N_XI42/XI520/XI16/NET048_XI42/XI520/XI16/MM18_d
+ N_NET136_XI42/XI520/XI16/MM18_g N_VSS_XI42/XI520/XI16/MM18_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13
+ AS=2.726e-13 PD=5.1e-07 PS=1.63e-06
mXI42/XI520/XI17/MM16 N_XI42/NET375_XI42/XI520/XI17/MM16_d
+ N_NET139_XI42/XI520/XI17/MM16_g
+ N_XI42/XI520/XI17/NET034_XI42/XI520/XI17/MM16_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI42/XI520/XI17/MM17 N_XI42/XI520/XI17/NET034_XI42/XI520/XI17/MM17_d
+ N_NET138_XI42/XI520/XI17/MM17_g
+ N_XI42/XI520/XI17/NET048_XI42/XI520/XI17/MM17_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13
+ AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI42/XI520/XI17/MM18 N_XI42/XI520/XI17/NET048_XI42/XI520/XI17/MM18_d
+ N_NET135_XI42/XI520/XI17/MM18_g N_VSS_XI42/XI520/XI17/MM18_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13
+ AS=2.726e-13 PD=5.1e-07 PS=1.63e-06
mXI42/XI520/XI18/MM16 N_XI42/NET535_XI42/XI520/XI18/MM16_d
+ N_NET139_XI42/XI520/XI18/MM16_g
+ N_XI42/XI520/XI18/NET034_XI42/XI520/XI18/MM16_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI42/XI520/XI18/MM17 N_XI42/XI520/XI18/NET034_XI42/XI520/XI18/MM17_d
+ N_NET137_XI42/XI520/XI18/MM17_g
+ N_XI42/XI520/XI18/NET048_XI42/XI520/XI18/MM17_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13
+ AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI42/XI520/XI18/MM18 N_XI42/XI520/XI18/NET048_XI42/XI520/XI18/MM18_d
+ N_NET136_XI42/XI520/XI18/MM18_g N_VSS_XI42/XI520/XI18/MM18_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13
+ AS=2.726e-13 PD=5.1e-07 PS=1.63e-06
mXI42/XI520/XI19/MM16 N_XI42/NET180_XI42/XI520/XI19/MM16_d
+ N_NET139_XI42/XI520/XI19/MM16_g
+ N_XI42/XI520/XI19/NET034_XI42/XI520/XI19/MM16_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI42/XI520/XI19/MM17 N_XI42/XI520/XI19/NET034_XI42/XI520/XI19/MM17_d
+ N_NET137_XI42/XI520/XI19/MM17_g
+ N_XI42/XI520/XI19/NET048_XI42/XI520/XI19/MM17_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13
+ AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI42/XI520/XI19/MM18 N_XI42/XI520/XI19/NET048_XI42/XI520/XI19/MM18_d
+ N_NET135_XI42/XI520/XI19/MM18_g N_VSS_XI42/XI520/XI19/MM18_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13
+ AS=2.726e-13 PD=5.1e-07 PS=1.63e-06
mXI54/XI0/XI8/XI3/MM2 N_XI54/XI0/XI8/NET12_XI54/XI0/XI8/XI3/MM2_d
+ N_NET068_XI54/XI0/XI8/XI3/MM2_g
+ N_XI54/XI0/XI8/XI3/NET13_XI54/XI0/XI8/XI3/MM2_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.3265e-13
+ AS=1.68025e-13 PD=1.46e-06 PS=7.15e-07
mXI54/XI0/XI7/XI3/MM2 N_XI54/XI0/XI7/NET12_XI54/XI0/XI7/XI3/MM2_d
+ N_NET068_XI54/XI0/XI7/XI3/MM2_g
+ N_XI54/XI0/XI7/XI3/NET13_XI54/XI0/XI7/XI3/MM2_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.3265e-13
+ AS=1.68025e-13 PD=1.46e-06 PS=7.15e-07
mXI54/XI0/XI8/XI3/MM3 N_XI54/XI0/XI8/XI3/NET13_XI54/XI0/XI8/XI3/MM3_d
+ N_XI54/XI0/NET2_XI54/XI0/XI8/XI3/MM3_g N_VSS_XI54/XI0/XI8/XI3/MM3_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=1.68025e-13
+ AS=2.303e-13 PD=7.15e-07 PS=1.45e-06
mXI54/XI0/XI7/XI3/MM3 N_XI54/XI0/XI7/XI3/NET13_XI54/XI0/XI7/XI3/MM3_d
+ N_NET062_XI54/XI0/XI7/XI3/MM3_g N_VSS_XI54/XI0/XI7/XI3/MM3_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=1.68025e-13
+ AS=2.303e-13 PD=7.15e-07 PS=1.45e-06
mXI54/XI0/XI6/MM1 N_XI54/XI0/NET2_XI54/XI0/XI6/MM1_d N_NET062_XI54/XI0/XI6/MM1_g
+ N_VSS_XI54/XI0/XI6/MM1_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI42/XI649/XI2/MM2 N_XI42/NET0373_XI42/XI649/XI2/MM2_d
+ N_NET070_XI42/XI649/XI2/MM2_g N_XI42/XI649/XI2/NET13_XI42/XI649/XI2/MM2_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.397e-13
+ AS=1.692e-13 PD=1.49e-06 PS=7.2e-07
mXI42/XI648/MM5 N_XI42/NET01023_XI42/XI648/MM5_d N_XI42/NET801_XI42/XI648/MM5_g
+ N_VSS_XI42/XI648/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI584/MM5 N_NET280_XI42/XI584/MM5_d N_XI42/NET455_XI42/XI584/MM5_g
+ N_VSS_XI42/XI584/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI616/MM5 N_NET281_XI42/XI616/MM5_d N_XI42/NET803_XI42/XI616/MM5_g
+ N_VSS_XI42/XI616/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI552/MM5 N_NET282_XI42/XI552/MM5_d N_XI42/NET245_XI42/XI552/MM5_g
+ N_VSS_XI42/XI552/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI632/MM5 N_NET153_XI42/XI632/MM5_d N_XI42/NET802_XI42/XI632/MM5_g
+ N_VSS_XI42/XI632/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI568/MM5 N_NET284_XI42/XI568/MM5_d N_XI42/NET375_XI42/XI568/MM5_g
+ N_VSS_XI42/XI568/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI600/MM5 N_NET285_XI42/XI600/MM5_d N_XI42/NET535_XI42/XI600/MM5_g
+ N_VSS_XI42/XI600/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI536/MM5 N_NET286_XI42/XI536/MM5_d N_XI42/NET180_XI42/XI536/MM5_g
+ N_VSS_XI42/XI536/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI647/MM5 N_NET287_XI42/XI647/MM5_d N_XI42/NET801_XI42/XI647/MM5_g
+ N_VSS_XI42/XI647/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI583/MM5 N_NET158_XI42/XI583/MM5_d N_XI42/NET455_XI42/XI583/MM5_g
+ N_VSS_XI42/XI583/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI615/MM5 N_NET159_XI42/XI615/MM5_d N_XI42/NET803_XI42/XI615/MM5_g
+ N_VSS_XI42/XI615/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI551/MM5 N_NET160_XI42/XI551/MM5_d N_XI42/NET245_XI42/XI551/MM5_g
+ N_VSS_XI42/XI551/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI631/MM5 N_NET291_XI42/XI631/MM5_d N_XI42/NET802_XI42/XI631/MM5_g
+ N_VSS_XI42/XI631/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI567/MM5 N_NET162_XI42/XI567/MM5_d N_XI42/NET375_XI42/XI567/MM5_g
+ N_VSS_XI42/XI567/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI599/MM5 N_NET293_XI42/XI599/MM5_d N_XI42/NET535_XI42/XI599/MM5_g
+ N_VSS_XI42/XI599/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI535/MM5 N_NET294_XI42/XI535/MM5_d N_XI42/NET180_XI42/XI535/MM5_g
+ N_VSS_XI42/XI535/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI646/MM5 N_NET295_XI42/XI646/MM5_d N_XI42/NET801_XI42/XI646/MM5_g
+ N_VSS_XI42/XI646/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI582/MM5 N_NET296_XI42/XI582/MM5_d N_XI42/NET455_XI42/XI582/MM5_g
+ N_VSS_XI42/XI582/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI614/MM5 N_NET297_XI42/XI614/MM5_d N_XI42/NET803_XI42/XI614/MM5_g
+ N_VSS_XI42/XI614/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI550/MM5 N_NET298_XI42/XI550/MM5_d N_XI42/NET245_XI42/XI550/MM5_g
+ N_VSS_XI42/XI550/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI630/MM5 N_NET299_XI42/XI630/MM5_d N_XI42/NET802_XI42/XI630/MM5_g
+ N_VSS_XI42/XI630/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI566/MM5 N_NET170_XI42/XI566/MM5_d N_XI42/NET375_XI42/XI566/MM5_g
+ N_VSS_XI42/XI566/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI598/MM5 N_NET171_XI42/XI598/MM5_d N_XI42/NET535_XI42/XI598/MM5_g
+ N_VSS_XI42/XI598/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI534/MM5 N_NET172_XI42/XI534/MM5_d N_XI42/NET180_XI42/XI534/MM5_g
+ N_VSS_XI42/XI534/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI645/MM5 N_NET303_XI42/XI645/MM5_d N_XI42/NET801_XI42/XI645/MM5_g
+ N_VSS_XI42/XI645/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI581/MM5 N_NET304_XI42/XI581/MM5_d N_XI42/NET455_XI42/XI581/MM5_g
+ N_VSS_XI42/XI581/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI613/MM5 N_NET305_XI42/XI613/MM5_d N_XI42/NET803_XI42/XI613/MM5_g
+ N_VSS_XI42/XI613/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI549/MM5 N_NET306_XI42/XI549/MM5_d N_XI42/NET245_XI42/XI549/MM5_g
+ N_VSS_XI42/XI549/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI629/MM5 N_NET307_XI42/XI629/MM5_d N_XI42/NET802_XI42/XI629/MM5_g
+ N_VSS_XI42/XI629/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI565/MM5 N_NET308_XI42/XI565/MM5_d N_XI42/NET375_XI42/XI565/MM5_g
+ N_VSS_XI42/XI565/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI597/MM5 N_NET309_XI42/XI597/MM5_d N_XI42/NET535_XI42/XI597/MM5_g
+ N_VSS_XI42/XI597/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI533/MM5 N_NET310_XI42/XI533/MM5_d N_XI42/NET180_XI42/XI533/MM5_g
+ N_VSS_XI42/XI533/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI644/MM5 N_NET311_XI42/XI644/MM5_d N_XI42/NET801_XI42/XI644/MM5_g
+ N_VSS_XI42/XI644/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI580/MM5 N_NET312_XI42/XI580/MM5_d N_XI42/NET455_XI42/XI580/MM5_g
+ N_VSS_XI42/XI580/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI612/MM5 N_NET313_XI42/XI612/MM5_d N_XI42/NET803_XI42/XI612/MM5_g
+ N_VSS_XI42/XI612/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI548/MM5 N_NET314_XI42/XI548/MM5_d N_XI42/NET245_XI42/XI548/MM5_g
+ N_VSS_XI42/XI548/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI628/MM5 N_NET315_XI42/XI628/MM5_d N_XI42/NET802_XI42/XI628/MM5_g
+ N_VSS_XI42/XI628/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI564/MM5 N_NET316_XI42/XI564/MM5_d N_XI42/NET375_XI42/XI564/MM5_g
+ N_VSS_XI42/XI564/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI596/MM5 N_NET317_XI42/XI596/MM5_d N_XI42/NET535_XI42/XI596/MM5_g
+ N_VSS_XI42/XI596/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI532/MM5 N_NET318_XI42/XI532/MM5_d N_XI42/NET180_XI42/XI532/MM5_g
+ N_VSS_XI42/XI532/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI643/MM5 N_NET319_XI42/XI643/MM5_d N_XI42/NET801_XI42/XI643/MM5_g
+ N_VSS_XI42/XI643/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI579/MM5 N_NET320_XI42/XI579/MM5_d N_XI42/NET455_XI42/XI579/MM5_g
+ N_VSS_XI42/XI579/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI611/MM5 N_NET321_XI42/XI611/MM5_d N_XI42/NET803_XI42/XI611/MM5_g
+ N_VSS_XI42/XI611/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI547/MM5 N_NET192_XI42/XI547/MM5_d N_XI42/NET245_XI42/XI547/MM5_g
+ N_VSS_XI42/XI547/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI627/MM5 N_NET193_XI42/XI627/MM5_d N_XI42/NET802_XI42/XI627/MM5_g
+ N_VSS_XI42/XI627/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI563/MM5 N_NET194_XI42/XI563/MM5_d N_XI42/NET375_XI42/XI563/MM5_g
+ N_VSS_XI42/XI563/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI595/MM5 N_NET195_XI42/XI595/MM5_d N_XI42/NET535_XI42/XI595/MM5_g
+ N_VSS_XI42/XI595/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI531/MM5 N_NET196_XI42/XI531/MM5_d N_XI42/NET180_XI42/XI531/MM5_g
+ N_VSS_XI42/XI531/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI642/MM5 N_NET197_XI42/XI642/MM5_d N_XI42/NET801_XI42/XI642/MM5_g
+ N_VSS_XI42/XI642/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI578/MM5 N_NET198_XI42/XI578/MM5_d N_XI42/NET455_XI42/XI578/MM5_g
+ N_VSS_XI42/XI578/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI610/MM5 N_NET199_XI42/XI610/MM5_d N_XI42/NET803_XI42/XI610/MM5_g
+ N_VSS_XI42/XI610/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI546/MM5 N_NET200_XI42/XI546/MM5_d N_XI42/NET245_XI42/XI546/MM5_g
+ N_VSS_XI42/XI546/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI626/MM5 N_NET331_XI42/XI626/MM5_d N_XI42/NET802_XI42/XI626/MM5_g
+ N_VSS_XI42/XI626/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI562/MM5 N_NET332_XI42/XI562/MM5_d N_XI42/NET375_XI42/XI562/MM5_g
+ N_VSS_XI42/XI562/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI594/MM5 N_NET203_XI42/XI594/MM5_d N_XI42/NET535_XI42/XI594/MM5_g
+ N_VSS_XI42/XI594/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI530/MM5 N_NET204_XI42/XI530/MM5_d N_XI42/NET180_XI42/XI530/MM5_g
+ N_VSS_XI42/XI530/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI641/MM5 N_NET205_XI42/XI641/MM5_d N_XI42/NET801_XI42/XI641/MM5_g
+ N_VSS_XI42/XI641/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI577/MM5 N_NET206_XI42/XI577/MM5_d N_XI42/NET455_XI42/XI577/MM5_g
+ N_VSS_XI42/XI577/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI609/MM5 N_NET207_XI42/XI609/MM5_d N_XI42/NET803_XI42/XI609/MM5_g
+ N_VSS_XI42/XI609/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI545/MM5 N_NET338_XI42/XI545/MM5_d N_XI42/NET245_XI42/XI545/MM5_g
+ N_VSS_XI42/XI545/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI625/MM5 N_NET339_XI42/XI625/MM5_d N_XI42/NET802_XI42/XI625/MM5_g
+ N_VSS_XI42/XI625/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI561/MM5 N_NET340_XI42/XI561/MM5_d N_XI42/NET375_XI42/XI561/MM5_g
+ N_VSS_XI42/XI561/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI593/MM5 N_NET211_XI42/XI593/MM5_d N_XI42/NET535_XI42/XI593/MM5_g
+ N_VSS_XI42/XI593/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI529/MM5 N_NET212_XI42/XI529/MM5_d N_XI42/NET180_XI42/XI529/MM5_g
+ N_VSS_XI42/XI529/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI640/MM5 N_NET214_XI42/XI640/MM5_d N_XI42/NET801_XI42/XI640/MM5_g
+ N_VSS_XI42/XI640/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI576/MM5 N_NET215_XI42/XI576/MM5_d N_XI42/NET455_XI42/XI576/MM5_g
+ N_VSS_XI42/XI576/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI608/MM5 N_NET216_XI42/XI608/MM5_d N_XI42/NET803_XI42/XI608/MM5_g
+ N_VSS_XI42/XI608/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI544/MM5 N_NET346_XI42/XI544/MM5_d N_XI42/NET245_XI42/XI544/MM5_g
+ N_VSS_XI42/XI544/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI624/MM5 N_NET347_XI42/XI624/MM5_d N_XI42/NET802_XI42/XI624/MM5_g
+ N_VSS_XI42/XI624/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI560/MM5 N_NET348_XI42/XI560/MM5_d N_XI42/NET375_XI42/XI560/MM5_g
+ N_VSS_XI42/XI560/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI592/MM5 N_NET349_XI42/XI592/MM5_d N_XI42/NET535_XI42/XI592/MM5_g
+ N_VSS_XI42/XI592/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI528/MM5 N_NET350_XI42/XI528/MM5_d N_XI42/NET180_XI42/XI528/MM5_g
+ N_VSS_XI42/XI528/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI639/MM5 N_NET351_XI42/XI639/MM5_d N_XI42/NET801_XI42/XI639/MM5_g
+ N_VSS_XI42/XI639/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI575/MM5 N_NET352_XI42/XI575/MM5_d N_XI42/NET455_XI42/XI575/MM5_g
+ N_VSS_XI42/XI575/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI607/MM5 N_NET224_XI42/XI607/MM5_d N_XI42/NET803_XI42/XI607/MM5_g
+ N_VSS_XI42/XI607/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI543/MM5 N_NET225_XI42/XI543/MM5_d N_XI42/NET245_XI42/XI543/MM5_g
+ N_VSS_XI42/XI543/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI623/MM5 N_NET226_XI42/XI623/MM5_d N_XI42/NET802_XI42/XI623/MM5_g
+ N_VSS_XI42/XI623/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI559/MM5 N_NET356_XI42/XI559/MM5_d N_XI42/NET375_XI42/XI559/MM5_g
+ N_VSS_XI42/XI559/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI591/MM5 N_NET357_XI42/XI591/MM5_d N_XI42/NET535_XI42/XI591/MM5_g
+ N_VSS_XI42/XI591/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI527/MM5 N_NET358_XI42/XI527/MM5_d N_XI42/NET180_XI42/XI527/MM5_g
+ N_VSS_XI42/XI527/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI638/MM5 N_NET230_XI42/XI638/MM5_d N_XI42/NET801_XI42/XI638/MM5_g
+ N_VSS_XI42/XI638/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI574/MM5 N_NET360_XI42/XI574/MM5_d N_XI42/NET455_XI42/XI574/MM5_g
+ N_VSS_XI42/XI574/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI606/MM5 N_NET361_XI42/XI606/MM5_d N_XI42/NET803_XI42/XI606/MM5_g
+ N_VSS_XI42/XI606/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI542/MM5 N_NET233_XI42/XI542/MM5_d N_XI42/NET245_XI42/XI542/MM5_g
+ N_VSS_XI42/XI542/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI622/MM5 N_NET234_XI42/XI622/MM5_d N_XI42/NET802_XI42/XI622/MM5_g
+ N_VSS_XI42/XI622/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI558/MM5 N_NET235_XI42/XI558/MM5_d N_XI42/NET375_XI42/XI558/MM5_g
+ N_VSS_XI42/XI558/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI590/MM5 N_NET365_XI42/XI590/MM5_d N_XI42/NET535_XI42/XI590/MM5_g
+ N_VSS_XI42/XI590/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI526/MM5 N_NET366_XI42/XI526/MM5_d N_XI42/NET180_XI42/XI526/MM5_g
+ N_VSS_XI42/XI526/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI637/MM5 N_NET367_XI42/XI637/MM5_d N_XI42/NET801_XI42/XI637/MM5_g
+ N_VSS_XI42/XI637/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI573/MM5 N_NET368_XI42/XI573/MM5_d N_XI42/NET455_XI42/XI573/MM5_g
+ N_VSS_XI42/XI573/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI605/MM5 N_NET369_XI42/XI605/MM5_d N_XI42/NET803_XI42/XI605/MM5_g
+ N_VSS_XI42/XI605/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI541/MM5 N_NET370_XI42/XI541/MM5_d N_XI42/NET245_XI42/XI541/MM5_g
+ N_VSS_XI42/XI541/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI621/MM5 N_NET371_XI42/XI621/MM5_d N_XI42/NET802_XI42/XI621/MM5_g
+ N_VSS_XI42/XI621/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI557/MM5 N_NET242_XI42/XI557/MM5_d N_XI42/NET375_XI42/XI557/MM5_g
+ N_VSS_XI42/XI557/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI589/MM5 N_NET373_XI42/XI589/MM5_d N_XI42/NET535_XI42/XI589/MM5_g
+ N_VSS_XI42/XI589/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI525/MM5 N_NET244_XI42/XI525/MM5_d N_XI42/NET180_XI42/XI525/MM5_g
+ N_VSS_XI42/XI525/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI636/MM5 N_NET375_XI42/XI636/MM5_d N_XI42/NET801_XI42/XI636/MM5_g
+ N_VSS_XI42/XI636/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI572/MM5 N_NET376_XI42/XI572/MM5_d N_XI42/NET455_XI42/XI572/MM5_g
+ N_VSS_XI42/XI572/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI604/MM5 N_NET377_XI42/XI604/MM5_d N_XI42/NET803_XI42/XI604/MM5_g
+ N_VSS_XI42/XI604/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI540/MM5 N_NET378_XI42/XI540/MM5_d N_XI42/NET245_XI42/XI540/MM5_g
+ N_VSS_XI42/XI540/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI620/MM5 N_NET379_XI42/XI620/MM5_d N_XI42/NET802_XI42/XI620/MM5_g
+ N_VSS_XI42/XI620/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI556/MM5 N_NET380_XI42/XI556/MM5_d N_XI42/NET375_XI42/XI556/MM5_g
+ N_VSS_XI42/XI556/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI588/MM5 N_NET381_XI42/XI588/MM5_d N_XI42/NET535_XI42/XI588/MM5_g
+ N_VSS_XI42/XI588/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI524/MM5 N_NET382_XI42/XI524/MM5_d N_XI42/NET180_XI42/XI524/MM5_g
+ N_VSS_XI42/XI524/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI635/MM5 N_NET383_XI42/XI635/MM5_d N_XI42/NET801_XI42/XI635/MM5_g
+ N_VSS_XI42/XI635/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI571/MM5 N_NET384_XI42/XI571/MM5_d N_XI42/NET455_XI42/XI571/MM5_g
+ N_VSS_XI42/XI571/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI603/MM5 N_NET385_XI42/XI603/MM5_d N_XI42/NET803_XI42/XI603/MM5_g
+ N_VSS_XI42/XI603/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI539/MM5 N_NET256_XI42/XI539/MM5_d N_XI42/NET245_XI42/XI539/MM5_g
+ N_VSS_XI42/XI539/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI619/MM5 N_NET387_XI42/XI619/MM5_d N_XI42/NET802_XI42/XI619/MM5_g
+ N_VSS_XI42/XI619/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI555/MM5 N_NET388_XI42/XI555/MM5_d N_XI42/NET375_XI42/XI555/MM5_g
+ N_VSS_XI42/XI555/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI587/MM5 N_NET389_XI42/XI587/MM5_d N_XI42/NET535_XI42/XI587/MM5_g
+ N_VSS_XI42/XI587/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI523/MM5 N_NET390_XI42/XI523/MM5_d N_XI42/NET180_XI42/XI523/MM5_g
+ N_VSS_XI42/XI523/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI634/MM5 N_NET391_XI42/XI634/MM5_d N_XI42/NET801_XI42/XI634/MM5_g
+ N_VSS_XI42/XI634/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI570/MM5 N_NET262_XI42/XI570/MM5_d N_XI42/NET455_XI42/XI570/MM5_g
+ N_VSS_XI42/XI570/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI602/MM5 N_NET263_XI42/XI602/MM5_d N_XI42/NET803_XI42/XI602/MM5_g
+ N_VSS_XI42/XI602/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI538/MM5 N_NET264_XI42/XI538/MM5_d N_XI42/NET245_XI42/XI538/MM5_g
+ N_VSS_XI42/XI538/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI618/MM5 N_NET265_XI42/XI618/MM5_d N_XI42/NET802_XI42/XI618/MM5_g
+ N_VSS_XI42/XI618/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI554/MM5 N_NET396_XI42/XI554/MM5_d N_XI42/NET375_XI42/XI554/MM5_g
+ N_VSS_XI42/XI554/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI586/MM5 N_NET267_XI42/XI586/MM5_d N_XI42/NET535_XI42/XI586/MM5_g
+ N_VSS_XI42/XI586/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI522/MM5 N_NET268_XI42/XI522/MM5_d N_XI42/NET180_XI42/XI522/MM5_g
+ N_VSS_XI42/XI522/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI633/MM5 N_NET269_XI42/XI633/MM5_d N_XI42/NET801_XI42/XI633/MM5_g
+ N_VSS_XI42/XI633/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI569/MM5 N_NET270_XI42/XI569/MM5_d N_XI42/NET455_XI42/XI569/MM5_g
+ N_VSS_XI42/XI569/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI601/MM5 N_NET401_XI42/XI601/MM5_d N_XI42/NET803_XI42/XI601/MM5_g
+ N_VSS_XI42/XI601/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI537/MM5 N_NET272_XI42/XI537/MM5_d N_XI42/NET245_XI42/XI537/MM5_g
+ N_VSS_XI42/XI537/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI617/MM5 N_NET273_XI42/XI617/MM5_d N_XI42/NET802_XI42/XI617/MM5_g
+ N_VSS_XI42/XI617/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI553/MM5 N_NET404_XI42/XI553/MM5_d N_XI42/NET375_XI42/XI553/MM5_g
+ N_VSS_XI42/XI553/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI585/MM5 N_NET405_XI42/XI585/MM5_d N_XI42/NET535_XI42/XI585/MM5_g
+ N_VSS_XI42/XI585/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI521/MM5 N_XI42/NET0388_XI42/XI521/MM5_d N_XI42/NET180_XI42/XI521/MM5_g
+ N_VSS_XI42/XI521/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI649/XI2/MM3 N_XI42/XI649/XI2/NET13_XI42/XI649/XI2/MM3_d
+ N_XI42/NET0388_XI42/XI649/XI2/MM3_g N_VSS_XI42/XI649/XI2/MM3_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13
+ AS=2.679e-13 PD=7.2e-07 PS=1.61e-06
mXI42/XI648/MM4 N_XI42/NET01023_XI42/XI648/MM4_d N_XI42/NET780_XI42/XI648/MM4_g
+ N_VSS_XI42/XI648/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI584/MM4 N_NET280_XI42/XI584/MM4_d N_XI42/NET780_XI42/XI584/MM4_g
+ N_VSS_XI42/XI584/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI616/MM4 N_NET281_XI42/XI616/MM4_d N_XI42/NET780_XI42/XI616/MM4_g
+ N_VSS_XI42/XI616/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI552/MM4 N_NET282_XI42/XI552/MM4_d N_XI42/NET780_XI42/XI552/MM4_g
+ N_VSS_XI42/XI552/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI632/MM4 N_NET153_XI42/XI632/MM4_d N_XI42/NET780_XI42/XI632/MM4_g
+ N_VSS_XI42/XI632/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI568/MM4 N_NET284_XI42/XI568/MM4_d N_XI42/NET780_XI42/XI568/MM4_g
+ N_VSS_XI42/XI568/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI600/MM4 N_NET285_XI42/XI600/MM4_d N_XI42/NET780_XI42/XI600/MM4_g
+ N_VSS_XI42/XI600/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI536/MM4 N_NET286_XI42/XI536/MM4_d N_XI42/NET780_XI42/XI536/MM4_g
+ N_VSS_XI42/XI536/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI647/MM4 N_NET287_XI42/XI647/MM4_d N_XI42/NET781_XI42/XI647/MM4_g
+ N_VSS_XI42/XI647/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI583/MM4 N_NET158_XI42/XI583/MM4_d N_XI42/NET781_XI42/XI583/MM4_g
+ N_VSS_XI42/XI583/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI615/MM4 N_NET159_XI42/XI615/MM4_d N_XI42/NET781_XI42/XI615/MM4_g
+ N_VSS_XI42/XI615/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI551/MM4 N_NET160_XI42/XI551/MM4_d N_XI42/NET781_XI42/XI551/MM4_g
+ N_VSS_XI42/XI551/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI631/MM4 N_NET291_XI42/XI631/MM4_d N_XI42/NET781_XI42/XI631/MM4_g
+ N_VSS_XI42/XI631/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI567/MM4 N_NET162_XI42/XI567/MM4_d N_XI42/NET781_XI42/XI567/MM4_g
+ N_VSS_XI42/XI567/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI599/MM4 N_NET293_XI42/XI599/MM4_d N_XI42/NET781_XI42/XI599/MM4_g
+ N_VSS_XI42/XI599/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI535/MM4 N_NET294_XI42/XI535/MM4_d N_XI42/NET781_XI42/XI535/MM4_g
+ N_VSS_XI42/XI535/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI646/MM4 N_NET295_XI42/XI646/MM4_d N_XI42/NET782_XI42/XI646/MM4_g
+ N_VSS_XI42/XI646/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI582/MM4 N_NET296_XI42/XI582/MM4_d N_XI42/NET782_XI42/XI582/MM4_g
+ N_VSS_XI42/XI582/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI614/MM4 N_NET297_XI42/XI614/MM4_d N_XI42/NET782_XI42/XI614/MM4_g
+ N_VSS_XI42/XI614/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI550/MM4 N_NET298_XI42/XI550/MM4_d N_XI42/NET782_XI42/XI550/MM4_g
+ N_VSS_XI42/XI550/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI630/MM4 N_NET299_XI42/XI630/MM4_d N_XI42/NET782_XI42/XI630/MM4_g
+ N_VSS_XI42/XI630/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI566/MM4 N_NET170_XI42/XI566/MM4_d N_XI42/NET782_XI42/XI566/MM4_g
+ N_VSS_XI42/XI566/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI598/MM4 N_NET171_XI42/XI598/MM4_d N_XI42/NET782_XI42/XI598/MM4_g
+ N_VSS_XI42/XI598/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI534/MM4 N_NET172_XI42/XI534/MM4_d N_XI42/NET782_XI42/XI534/MM4_g
+ N_VSS_XI42/XI534/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI645/MM4 N_NET303_XI42/XI645/MM4_d N_XI42/NET783_XI42/XI645/MM4_g
+ N_VSS_XI42/XI645/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI581/MM4 N_NET304_XI42/XI581/MM4_d N_XI42/NET783_XI42/XI581/MM4_g
+ N_VSS_XI42/XI581/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI613/MM4 N_NET305_XI42/XI613/MM4_d N_XI42/NET783_XI42/XI613/MM4_g
+ N_VSS_XI42/XI613/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI549/MM4 N_NET306_XI42/XI549/MM4_d N_XI42/NET783_XI42/XI549/MM4_g
+ N_VSS_XI42/XI549/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI629/MM4 N_NET307_XI42/XI629/MM4_d N_XI42/NET783_XI42/XI629/MM4_g
+ N_VSS_XI42/XI629/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI565/MM4 N_NET308_XI42/XI565/MM4_d N_XI42/NET783_XI42/XI565/MM4_g
+ N_VSS_XI42/XI565/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI597/MM4 N_NET309_XI42/XI597/MM4_d N_XI42/NET783_XI42/XI597/MM4_g
+ N_VSS_XI42/XI597/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI533/MM4 N_NET310_XI42/XI533/MM4_d N_XI42/NET783_XI42/XI533/MM4_g
+ N_VSS_XI42/XI533/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI644/MM4 N_NET311_XI42/XI644/MM4_d N_XI42/NET784_XI42/XI644/MM4_g
+ N_VSS_XI42/XI644/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI580/MM4 N_NET312_XI42/XI580/MM4_d N_XI42/NET784_XI42/XI580/MM4_g
+ N_VSS_XI42/XI580/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI612/MM4 N_NET313_XI42/XI612/MM4_d N_XI42/NET784_XI42/XI612/MM4_g
+ N_VSS_XI42/XI612/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI548/MM4 N_NET314_XI42/XI548/MM4_d N_XI42/NET784_XI42/XI548/MM4_g
+ N_VSS_XI42/XI548/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI628/MM4 N_NET315_XI42/XI628/MM4_d N_XI42/NET784_XI42/XI628/MM4_g
+ N_VSS_XI42/XI628/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI564/MM4 N_NET316_XI42/XI564/MM4_d N_XI42/NET784_XI42/XI564/MM4_g
+ N_VSS_XI42/XI564/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI596/MM4 N_NET317_XI42/XI596/MM4_d N_XI42/NET784_XI42/XI596/MM4_g
+ N_VSS_XI42/XI596/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI532/MM4 N_NET318_XI42/XI532/MM4_d N_XI42/NET784_XI42/XI532/MM4_g
+ N_VSS_XI42/XI532/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI643/MM4 N_NET319_XI42/XI643/MM4_d N_XI42/NET785_XI42/XI643/MM4_g
+ N_VSS_XI42/XI643/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI579/MM4 N_NET320_XI42/XI579/MM4_d N_XI42/NET785_XI42/XI579/MM4_g
+ N_VSS_XI42/XI579/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI611/MM4 N_NET321_XI42/XI611/MM4_d N_XI42/NET785_XI42/XI611/MM4_g
+ N_VSS_XI42/XI611/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI547/MM4 N_NET192_XI42/XI547/MM4_d N_XI42/NET785_XI42/XI547/MM4_g
+ N_VSS_XI42/XI547/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI627/MM4 N_NET193_XI42/XI627/MM4_d N_XI42/NET785_XI42/XI627/MM4_g
+ N_VSS_XI42/XI627/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI563/MM4 N_NET194_XI42/XI563/MM4_d N_XI42/NET785_XI42/XI563/MM4_g
+ N_VSS_XI42/XI563/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI595/MM4 N_NET195_XI42/XI595/MM4_d N_XI42/NET785_XI42/XI595/MM4_g
+ N_VSS_XI42/XI595/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI531/MM4 N_NET196_XI42/XI531/MM4_d N_XI42/NET785_XI42/XI531/MM4_g
+ N_VSS_XI42/XI531/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI642/MM4 N_NET197_XI42/XI642/MM4_d N_XI42/NET786_XI42/XI642/MM4_g
+ N_VSS_XI42/XI642/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI578/MM4 N_NET198_XI42/XI578/MM4_d N_XI42/NET786_XI42/XI578/MM4_g
+ N_VSS_XI42/XI578/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI610/MM4 N_NET199_XI42/XI610/MM4_d N_XI42/NET786_XI42/XI610/MM4_g
+ N_VSS_XI42/XI610/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI546/MM4 N_NET200_XI42/XI546/MM4_d N_XI42/NET786_XI42/XI546/MM4_g
+ N_VSS_XI42/XI546/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI626/MM4 N_NET331_XI42/XI626/MM4_d N_XI42/NET786_XI42/XI626/MM4_g
+ N_VSS_XI42/XI626/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI562/MM4 N_NET332_XI42/XI562/MM4_d N_XI42/NET786_XI42/XI562/MM4_g
+ N_VSS_XI42/XI562/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI594/MM4 N_NET203_XI42/XI594/MM4_d N_XI42/NET786_XI42/XI594/MM4_g
+ N_VSS_XI42/XI594/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI530/MM4 N_NET204_XI42/XI530/MM4_d N_XI42/NET786_XI42/XI530/MM4_g
+ N_VSS_XI42/XI530/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI641/MM4 N_NET205_XI42/XI641/MM4_d N_XI42/NET787_XI42/XI641/MM4_g
+ N_VSS_XI42/XI641/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI577/MM4 N_NET206_XI42/XI577/MM4_d N_XI42/NET787_XI42/XI577/MM4_g
+ N_VSS_XI42/XI577/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI609/MM4 N_NET207_XI42/XI609/MM4_d N_XI42/NET787_XI42/XI609/MM4_g
+ N_VSS_XI42/XI609/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI545/MM4 N_NET338_XI42/XI545/MM4_d N_XI42/NET787_XI42/XI545/MM4_g
+ N_VSS_XI42/XI545/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI625/MM4 N_NET339_XI42/XI625/MM4_d N_XI42/NET787_XI42/XI625/MM4_g
+ N_VSS_XI42/XI625/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI561/MM4 N_NET340_XI42/XI561/MM4_d N_XI42/NET787_XI42/XI561/MM4_g
+ N_VSS_XI42/XI561/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI593/MM4 N_NET211_XI42/XI593/MM4_d N_XI42/NET787_XI42/XI593/MM4_g
+ N_VSS_XI42/XI593/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI529/MM4 N_NET212_XI42/XI529/MM4_d N_XI42/NET787_XI42/XI529/MM4_g
+ N_VSS_XI42/XI529/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI640/MM4 N_NET214_XI42/XI640/MM4_d N_XI42/NET788_XI42/XI640/MM4_g
+ N_VSS_XI42/XI640/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI576/MM4 N_NET215_XI42/XI576/MM4_d N_XI42/NET788_XI42/XI576/MM4_g
+ N_VSS_XI42/XI576/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI608/MM4 N_NET216_XI42/XI608/MM4_d N_XI42/NET788_XI42/XI608/MM4_g
+ N_VSS_XI42/XI608/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI544/MM4 N_NET346_XI42/XI544/MM4_d N_XI42/NET788_XI42/XI544/MM4_g
+ N_VSS_XI42/XI544/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI624/MM4 N_NET347_XI42/XI624/MM4_d N_XI42/NET788_XI42/XI624/MM4_g
+ N_VSS_XI42/XI624/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI560/MM4 N_NET348_XI42/XI560/MM4_d N_XI42/NET788_XI42/XI560/MM4_g
+ N_VSS_XI42/XI560/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI592/MM4 N_NET349_XI42/XI592/MM4_d N_XI42/NET788_XI42/XI592/MM4_g
+ N_VSS_XI42/XI592/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI528/MM4 N_NET350_XI42/XI528/MM4_d N_XI42/NET788_XI42/XI528/MM4_g
+ N_VSS_XI42/XI528/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI639/MM4 N_NET351_XI42/XI639/MM4_d N_XI42/NET789_XI42/XI639/MM4_g
+ N_VSS_XI42/XI639/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI575/MM4 N_NET352_XI42/XI575/MM4_d N_XI42/NET789_XI42/XI575/MM4_g
+ N_VSS_XI42/XI575/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI607/MM4 N_NET224_XI42/XI607/MM4_d N_XI42/NET789_XI42/XI607/MM4_g
+ N_VSS_XI42/XI607/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI543/MM4 N_NET225_XI42/XI543/MM4_d N_XI42/NET789_XI42/XI543/MM4_g
+ N_VSS_XI42/XI543/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI623/MM4 N_NET226_XI42/XI623/MM4_d N_XI42/NET789_XI42/XI623/MM4_g
+ N_VSS_XI42/XI623/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI559/MM4 N_NET356_XI42/XI559/MM4_d N_XI42/NET789_XI42/XI559/MM4_g
+ N_VSS_XI42/XI559/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI591/MM4 N_NET357_XI42/XI591/MM4_d N_XI42/NET789_XI42/XI591/MM4_g
+ N_VSS_XI42/XI591/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI527/MM4 N_NET358_XI42/XI527/MM4_d N_XI42/NET789_XI42/XI527/MM4_g
+ N_VSS_XI42/XI527/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI638/MM4 N_NET230_XI42/XI638/MM4_d N_XI42/NET790_XI42/XI638/MM4_g
+ N_VSS_XI42/XI638/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI574/MM4 N_NET360_XI42/XI574/MM4_d N_XI42/NET790_XI42/XI574/MM4_g
+ N_VSS_XI42/XI574/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI606/MM4 N_NET361_XI42/XI606/MM4_d N_XI42/NET790_XI42/XI606/MM4_g
+ N_VSS_XI42/XI606/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI542/MM4 N_NET233_XI42/XI542/MM4_d N_XI42/NET790_XI42/XI542/MM4_g
+ N_VSS_XI42/XI542/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI622/MM4 N_NET234_XI42/XI622/MM4_d N_XI42/NET790_XI42/XI622/MM4_g
+ N_VSS_XI42/XI622/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI558/MM4 N_NET235_XI42/XI558/MM4_d N_XI42/NET790_XI42/XI558/MM4_g
+ N_VSS_XI42/XI558/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI590/MM4 N_NET365_XI42/XI590/MM4_d N_XI42/NET790_XI42/XI590/MM4_g
+ N_VSS_XI42/XI590/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI526/MM4 N_NET366_XI42/XI526/MM4_d N_XI42/NET790_XI42/XI526/MM4_g
+ N_VSS_XI42/XI526/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI637/MM4 N_NET367_XI42/XI637/MM4_d N_XI42/NET791_XI42/XI637/MM4_g
+ N_VSS_XI42/XI637/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI573/MM4 N_NET368_XI42/XI573/MM4_d N_XI42/NET791_XI42/XI573/MM4_g
+ N_VSS_XI42/XI573/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI605/MM4 N_NET369_XI42/XI605/MM4_d N_XI42/NET791_XI42/XI605/MM4_g
+ N_VSS_XI42/XI605/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI541/MM4 N_NET370_XI42/XI541/MM4_d N_XI42/NET791_XI42/XI541/MM4_g
+ N_VSS_XI42/XI541/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI621/MM4 N_NET371_XI42/XI621/MM4_d N_XI42/NET791_XI42/XI621/MM4_g
+ N_VSS_XI42/XI621/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI557/MM4 N_NET242_XI42/XI557/MM4_d N_XI42/NET791_XI42/XI557/MM4_g
+ N_VSS_XI42/XI557/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI589/MM4 N_NET373_XI42/XI589/MM4_d N_XI42/NET791_XI42/XI589/MM4_g
+ N_VSS_XI42/XI589/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI525/MM4 N_NET244_XI42/XI525/MM4_d N_XI42/NET791_XI42/XI525/MM4_g
+ N_VSS_XI42/XI525/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI636/MM4 N_NET375_XI42/XI636/MM4_d N_XI42/NET792_XI42/XI636/MM4_g
+ N_VSS_XI42/XI636/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI572/MM4 N_NET376_XI42/XI572/MM4_d N_XI42/NET792_XI42/XI572/MM4_g
+ N_VSS_XI42/XI572/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI604/MM4 N_NET377_XI42/XI604/MM4_d N_XI42/NET792_XI42/XI604/MM4_g
+ N_VSS_XI42/XI604/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI540/MM4 N_NET378_XI42/XI540/MM4_d N_XI42/NET792_XI42/XI540/MM4_g
+ N_VSS_XI42/XI540/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI620/MM4 N_NET379_XI42/XI620/MM4_d N_XI42/NET792_XI42/XI620/MM4_g
+ N_VSS_XI42/XI620/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI556/MM4 N_NET380_XI42/XI556/MM4_d N_XI42/NET792_XI42/XI556/MM4_g
+ N_VSS_XI42/XI556/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI588/MM4 N_NET381_XI42/XI588/MM4_d N_XI42/NET792_XI42/XI588/MM4_g
+ N_VSS_XI42/XI588/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI524/MM4 N_NET382_XI42/XI524/MM4_d N_XI42/NET792_XI42/XI524/MM4_g
+ N_VSS_XI42/XI524/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI635/MM4 N_NET383_XI42/XI635/MM4_d N_XI42/NET793_XI42/XI635/MM4_g
+ N_VSS_XI42/XI635/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI571/MM4 N_NET384_XI42/XI571/MM4_d N_XI42/NET793_XI42/XI571/MM4_g
+ N_VSS_XI42/XI571/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI603/MM4 N_NET385_XI42/XI603/MM4_d N_XI42/NET793_XI42/XI603/MM4_g
+ N_VSS_XI42/XI603/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI539/MM4 N_NET256_XI42/XI539/MM4_d N_XI42/NET793_XI42/XI539/MM4_g
+ N_VSS_XI42/XI539/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI619/MM4 N_NET387_XI42/XI619/MM4_d N_XI42/NET793_XI42/XI619/MM4_g
+ N_VSS_XI42/XI619/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI555/MM4 N_NET388_XI42/XI555/MM4_d N_XI42/NET793_XI42/XI555/MM4_g
+ N_VSS_XI42/XI555/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI587/MM4 N_NET389_XI42/XI587/MM4_d N_XI42/NET793_XI42/XI587/MM4_g
+ N_VSS_XI42/XI587/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI523/MM4 N_NET390_XI42/XI523/MM4_d N_XI42/NET793_XI42/XI523/MM4_g
+ N_VSS_XI42/XI523/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI634/MM4 N_NET391_XI42/XI634/MM4_d N_XI42/NET794_XI42/XI634/MM4_g
+ N_VSS_XI42/XI634/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI570/MM4 N_NET262_XI42/XI570/MM4_d N_XI42/NET794_XI42/XI570/MM4_g
+ N_VSS_XI42/XI570/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI602/MM4 N_NET263_XI42/XI602/MM4_d N_XI42/NET794_XI42/XI602/MM4_g
+ N_VSS_XI42/XI602/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI538/MM4 N_NET264_XI42/XI538/MM4_d N_XI42/NET794_XI42/XI538/MM4_g
+ N_VSS_XI42/XI538/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI618/MM4 N_NET265_XI42/XI618/MM4_d N_XI42/NET794_XI42/XI618/MM4_g
+ N_VSS_XI42/XI618/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI554/MM4 N_NET396_XI42/XI554/MM4_d N_XI42/NET794_XI42/XI554/MM4_g
+ N_VSS_XI42/XI554/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI586/MM4 N_NET267_XI42/XI586/MM4_d N_XI42/NET794_XI42/XI586/MM4_g
+ N_VSS_XI42/XI586/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI522/MM4 N_NET268_XI42/XI522/MM4_d N_XI42/NET794_XI42/XI522/MM4_g
+ N_VSS_XI42/XI522/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI633/MM4 N_NET269_XI42/XI633/MM4_d N_XI42/NET795_XI42/XI633/MM4_g
+ N_VSS_XI42/XI633/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI569/MM4 N_NET270_XI42/XI569/MM4_d N_XI42/NET795_XI42/XI569/MM4_g
+ N_VSS_XI42/XI569/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI601/MM4 N_NET401_XI42/XI601/MM4_d N_XI42/NET795_XI42/XI601/MM4_g
+ N_VSS_XI42/XI601/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI537/MM4 N_NET272_XI42/XI537/MM4_d N_XI42/NET795_XI42/XI537/MM4_g
+ N_VSS_XI42/XI537/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI617/MM4 N_NET273_XI42/XI617/MM4_d N_XI42/NET795_XI42/XI617/MM4_g
+ N_VSS_XI42/XI617/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI553/MM4 N_NET404_XI42/XI553/MM4_d N_XI42/NET795_XI42/XI553/MM4_g
+ N_VSS_XI42/XI553/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI585/MM4 N_NET405_XI42/XI585/MM4_d N_XI42/NET795_XI42/XI585/MM4_g
+ N_VSS_XI42/XI585/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI42/XI521/MM4 N_XI42/NET0388_XI42/XI521/MM4_d N_XI42/NET795_XI42/XI521/MM4_g
+ N_VSS_XI42/XI521/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.269e-13 AS=2.397e-13 PD=5.4e-07 PS=1.49e-06
mXI57/XI0/MM7 N_XI57/XI0/NET1_XI57/XI0/MM7_d N_NET064_XI57/XI0/MM7_g
+ N_XI57/XI0/NET9_XI57/XI0/MM7_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=1.2e-06 AD=4.5e-13 AS=6e-13 PD=7.5e-07 PS=2.2e-06
mXI57/XI0/MM5 N_XI57/NET19_XI57/XI0/MM5_d N_NET062_XI57/XI0/MM5_g
+ N_XI57/XI0/NET1_XI57/XI0/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=1.2e-06 AD=6.06e-13 AS=4.5e-13 PD=2.21e-06 PS=7.5e-07
mXI57/XI0/MM4 N_NET062_XI57/XI0/MM4_d N_XI57/NET19_XI57/XI0/MM4_g
+ N_XI57/XI0/NET20_XI57/XI0/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18
+ L=1.8e-07 W=1.2e-06 AD=6.06e-13 AS=4.5e-13 PD=2.21e-06 PS=7.5e-07
mXI57/XI0/MM6 N_XI57/XI0/NET20_XI57/XI0/MM6_d N_VREF_XI57/XI0/MM6_g
+ N_XI57/XI0/NET9_XI57/XI0/MM6_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=1.2e-06 AD=4.5e-13 AS=6e-13 PD=7.5e-07 PS=2.2e-06
mXI42/XI649/XI3/MM1 N_NET0390_XI42/XI649/XI3/MM1_d
+ N_XI42/NET0373_XI42/XI649/XI3/MM1_g N_VSS_XI42/XI649/XI3/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13
+ AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI57/XI0/MM8 N_XI57/XI0/NET9_XI57/XI0/MM8_d N_NET068_XI57/XI0/MM8_g
+ N_VSS_XI57/XI0/MM8_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI39/MM4095 N_NET0380_XI39/MM4095_d N_NET0133_XI39/MM4095_g N_VSS_XI39/MM4095_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3393 XI39/NET5650 N_NET280_XI39/MM3393_g N_VSS_XI39/MM3393_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3438 N_NET0380_XI39/MM3438_d N_NET281_XI39/MM3438_g N_VSS_XI39/MM3438_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3439 XI39/NET5466 N_NET282_XI39/MM3439_g N_VSS_XI39/MM3439_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3375 N_NET0380_XI39/MM3375_d N_NET153_XI39/MM3375_g N_VSS_XI39/MM3375_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3376 XI39/NET5718 N_NET284_XI39/MM3376_g N_VSS_XI39/MM3376_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3344 N_NET0380_XI39/MM3344_d N_NET285_XI39/MM3344_g N_VSS_XI39/MM3344_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3337 XI39/NET3574 N_NET286_XI39/MM3337_g N_VSS_XI39/MM3337_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3502 N_NET0380_XI39/MM3502_d N_NET287_XI39/MM3502_g N_VSS_XI39/MM3502_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3503 XI39/NET5210 N_NET158_XI39/MM3503_g N_VSS_XI39/MM3503_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3471 N_NET0380_XI39/MM3471_d N_NET159_XI39/MM3471_g N_VSS_XI39/MM3471_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3456 XI39/NET5398 N_NET160_XI39/MM3456_g N_VSS_XI39/MM3456_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3535 N_NET0380_XI39/MM3535_d N_NET291_XI39/MM3535_g N_VSS_XI39/MM3535_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3520 XI39/NET5142 N_NET162_XI39/MM3520_g N_VSS_XI39/MM3520_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3566 N_NET0380_XI39/MM3566_d N_NET293_XI39/MM3566_g N_VSS_XI39/MM3566_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3567 XI39/NET4954 N_NET294_XI39/MM3567_g N_VSS_XI39/MM3567_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3247 N_NET0380_XI39/MM3247_d N_NET295_XI39/MM3247_g N_VSS_XI39/MM3247_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3248 XI39/NET3930 N_NET296_XI39/MM3248_g N_VSS_XI39/MM3248_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3216 N_NET0380_XI39/MM3216_d N_NET297_XI39/MM3216_g N_VSS_XI39/MM3216_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3201 XI39/NET4118 N_NET298_XI39/MM3201_g N_VSS_XI39/MM3201_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3280 N_NET0380_XI39/MM3280_d N_NET299_XI39/MM3280_g N_VSS_XI39/MM3280_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3265 XI39/NET3862 N_NET170_XI39/MM3265_g N_VSS_XI39/MM3265_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3311 N_NET0380_XI39/MM3311_d N_NET171_XI39/MM3311_g N_VSS_XI39/MM3311_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3312 XI39/NET3674 N_NET172_XI39/MM3312_g N_VSS_XI39/MM3312_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3152 N_NET0380_XI39/MM3152_d N_NET303_XI39/MM3152_g N_VSS_XI39/MM3152_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3137 XI39/NET4374 N_NET304_XI39/MM3137_g N_VSS_XI39/MM3137_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3183 N_NET0380_XI39/MM3183_d N_NET305_XI39/MM3183_g N_VSS_XI39/MM3183_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3184 XI39/NET4186 N_NET306_XI39/MM3184_g N_VSS_XI39/MM3184_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3119 N_NET0380_XI39/MM3119_d N_NET307_XI39/MM3119_g N_VSS_XI39/MM3119_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3120 XI39/NET4442 N_NET308_XI39/MM3120_g N_VSS_XI39/MM3120_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3088 N_NET0380_XI39/MM3088_d N_NET309_XI39/MM3088_g N_VSS_XI39/MM3088_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3073 XI39/NET4630 N_NET310_XI39/MM3073_g N_VSS_XI39/MM3073_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3848 N_NET0380_XI39/MM3848_d N_NET311_XI39/MM3848_g N_VSS_XI39/MM3848_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3849 XI39/NET6126 N_NET312_XI39/MM3849_g N_VSS_XI39/MM3849_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3979 N_NET0380_XI39/MM3979_d N_NET313_XI39/MM3979_g N_VSS_XI39/MM3979_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3964 XI39/NET7462 N_NET314_XI39/MM3964_g N_VSS_XI39/MM3964_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3881 N_NET0380_XI39/MM3881_d N_NET315_XI39/MM3881_g N_VSS_XI39/MM3881_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3866 XI39/NET6058 N_NET316_XI39/MM3866_g N_VSS_XI39/MM3866_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3912 N_NET0380_XI39/MM3912_d N_NET317_XI39/MM3912_g N_VSS_XI39/MM3912_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3913 XI39/NET5870 N_NET318_XI39/MM3913_g N_VSS_XI39/MM3913_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4059 N_NET0380_XI39/MM4059_d N_NET319_XI39/MM4059_g N_VSS_XI39/MM4059_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4044 XI39/NET7142 N_NET320_XI39/MM4044_g N_VSS_XI39/MM4044_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3946 N_NET0380_XI39/MM3946_d N_NET321_XI39/MM3946_g N_VSS_XI39/MM3946_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3947 XI39/NET7530 N_NET192_XI39/MM3947_g N_VSS_XI39/MM3947_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4026 N_NET0380_XI39/MM4026_d N_NET193_XI39/MM4026_g N_VSS_XI39/MM4026_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4027 XI39/NET7210 N_NET194_XI39/MM4027_g N_VSS_XI39/MM4027_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4089 N_NET0380_XI39/MM4089_d N_NET195_XI39/MM4089_g N_VSS_XI39/MM4089_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4074 XI39/NET7022 N_NET196_XI39/MM4074_g N_VSS_XI39/MM4074_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3791 N_NET0380_XI39/MM3791_d N_NET197_XI39/MM3791_g N_VSS_XI39/MM3791_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3776 XI39/NET6418 N_NET198_XI39/MM3776_g N_VSS_XI39/MM3776_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3822 N_NET0380_XI39/MM3822_d N_NET199_XI39/MM3822_g N_VSS_XI39/MM3822_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3823 XI39/NET6230 N_NET200_XI39/MM3823_g N_VSS_XI39/MM3823_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3758 N_NET0380_XI39/MM3758_d N_NET331_XI39/MM3758_g N_VSS_XI39/MM3758_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3759 XI39/NET6486 N_NET332_XI39/MM3759_g N_VSS_XI39/MM3759_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3727 N_NET0380_XI39/MM3727_d N_NET203_XI39/MM3727_g N_VSS_XI39/MM3727_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3712 XI39/NET6674 N_NET204_XI39/MM3712_g N_VSS_XI39/MM3712_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3630 N_NET0380_XI39/MM3630_d N_NET205_XI39/MM3630_g N_VSS_XI39/MM3630_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3631 XI39/NET4698 N_NET206_XI39/MM3631_g N_VSS_XI39/MM3631_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3599 N_NET0380_XI39/MM3599_d N_NET207_XI39/MM3599_g N_VSS_XI39/MM3599_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3584 XI39/NET4886 N_NET338_XI39/MM3584_g N_VSS_XI39/MM3584_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3663 N_NET0380_XI39/MM3663_d N_NET339_XI39/MM3663_g N_VSS_XI39/MM3663_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3648 XI39/NET6930 N_NET340_XI39/MM3648_g N_VSS_XI39/MM3648_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3679 N_NET0380_XI39/MM3679_d N_NET211_XI39/MM3679_g N_VSS_XI39/MM3679_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3688 XI39/NET6770 N_NET212_XI39/MM3688_g N_VSS_XI39/MM3688_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2735 N_NET0380_XI39/MM2735_d N_NET214_XI39/MM2735_g N_VSS_XI39/MM2735_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2736 XI39/NET8922 N_NET215_XI39/MM2736_g N_VSS_XI39/MM2736_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2704 N_NET0380_XI39/MM2704_d N_NET216_XI39/MM2704_g N_VSS_XI39/MM2704_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2689 XI39/NET9106 N_NET346_XI39/MM2689_g N_VSS_XI39/MM2689_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2768 N_NET0380_XI39/MM2768_d N_NET347_XI39/MM2768_g N_VSS_XI39/MM2768_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2753 XI39/NET8854 N_NET348_XI39/MM2753_g N_VSS_XI39/MM2753_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2799 N_NET0380_XI39/MM2799_d N_NET349_XI39/MM2799_g N_VSS_XI39/MM2799_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2800 XI39/NET8666 N_NET350_XI39/MM2800_g N_VSS_XI39/MM2800_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2640 N_NET0380_XI39/MM2640_d N_NET351_XI39/MM2640_g N_VSS_XI39/MM2640_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2625 XI39/NET9362 N_NET352_XI39/MM2625_g N_VSS_XI39/MM2625_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2671 N_NET0380_XI39/MM2671_d N_NET224_XI39/MM2671_g N_VSS_XI39/MM2671_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2672 XI39/NET9174 N_NET225_XI39/MM2672_g N_VSS_XI39/MM2672_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2607 N_NET0380_XI39/MM2607_d N_NET226_XI39/MM2607_g N_VSS_XI39/MM2607_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2608 XI39/NET9430 N_NET356_XI39/MM2608_g N_VSS_XI39/MM2608_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2576 N_NET0380_XI39/MM2576_d N_NET357_XI39/MM2576_g N_VSS_XI39/MM2576_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2561 XI39/NET9618 N_NET358_XI39/MM2561_g N_VSS_XI39/MM2561_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2896 N_NET0380_XI39/MM2896_d N_NET230_XI39/MM2896_g N_VSS_XI39/MM2896_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2881 XI39/NET8342 N_NET360_XI39/MM2881_g N_VSS_XI39/MM2881_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2927 N_NET0380_XI39/MM2927_d N_NET361_XI39/MM2927_g N_VSS_XI39/MM2927_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2928 XI39/NET8154 N_NET233_XI39/MM2928_g N_VSS_XI39/MM2928_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2863 N_NET0380_XI39/MM2863_d N_NET234_XI39/MM2863_g N_VSS_XI39/MM2863_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2864 XI39/NET8410 N_NET235_XI39/MM2864_g N_VSS_XI39/MM2864_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2832 N_NET0380_XI39/MM2832_d N_NET365_XI39/MM2832_g N_VSS_XI39/MM2832_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2817 XI39/NET8598 N_NET366_XI39/MM2817_g N_VSS_XI39/MM2817_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2991 N_NET0380_XI39/MM2991_d N_NET367_XI39/MM2991_g N_VSS_XI39/MM2991_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2992 XI39/NET7898 N_NET368_XI39/MM2992_g N_VSS_XI39/MM2992_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2960 N_NET0380_XI39/MM2960_d N_NET369_XI39/MM2960_g N_VSS_XI39/MM2960_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2945 XI39/NET8086 N_NET370_XI39/MM2945_g N_VSS_XI39/MM2945_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3024 N_NET0380_XI39/MM3024_d N_NET371_XI39/MM3024_g N_VSS_XI39/MM3024_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3009 XI39/NET7830 N_NET242_XI39/MM3009_g N_VSS_XI39/MM3009_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3055 N_NET0380_XI39/MM3055_d N_NET373_XI39/MM3055_g N_VSS_XI39/MM3055_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3056 XI39/NET7642 N_NET244_XI39/MM3056_g N_VSS_XI39/MM3056_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2384 N_NET0380_XI39/MM2384_d N_NET375_XI39/MM2384_g N_VSS_XI39/MM2384_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2369 XI39/NET10746 N_NET376_XI39/MM2369_g N_VSS_XI39/MM2369_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2415 N_NET0380_XI39/MM2415_d N_NET377_XI39/MM2415_g N_VSS_XI39/MM2415_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2416 XI39/NET11206 N_NET378_XI39/MM2416_g N_VSS_XI39/MM2416_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2351 N_NET0380_XI39/MM2351_d N_NET379_XI39/MM2351_g N_VSS_XI39/MM2351_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2352 XI39/NET10814 N_NET380_XI39/MM2352_g N_VSS_XI39/MM2352_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2320 N_NET0380_XI39/MM2320_d N_NET381_XI39/MM2320_g N_VSS_XI39/MM2320_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2305 XI39/NET11002 N_NET382_XI39/MM2305_g N_VSS_XI39/MM2305_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2479 N_NET0380_XI39/MM2479_d N_NET383_XI39/MM2479_g N_VSS_XI39/MM2479_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2480 XI39/NET11526 N_NET384_XI39/MM2480_g N_VSS_XI39/MM2480_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2448 N_NET0380_XI39/MM2448_d N_NET385_XI39/MM2448_g N_VSS_XI39/MM2448_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2433 XI39/NET11138 N_NET256_XI39/MM2433_g N_VSS_XI39/MM2433_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2512 N_NET0380_XI39/MM2512_d N_NET387_XI39/MM2512_g N_VSS_XI39/MM2512_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2497 XI39/NET11458 N_NET388_XI39/MM2497_g N_VSS_XI39/MM2497_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2543 N_NET0380_XI39/MM2543_d N_NET389_XI39/MM2543_g N_VSS_XI39/MM2543_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2544 XI39/NET11646 N_NET390_XI39/MM2544_g N_VSS_XI39/MM2544_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4103 N_NET0380_XI39/MM4103_d N_NET391_XI39/MM4103_g N_VSS_XI39/MM4103_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2224 XI39/NET10458 N_NET262_XI39/MM2224_g N_VSS_XI39/MM2224_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4097 N_NET0380_XI39/MM4097_d N_NET263_XI39/MM4097_g N_VSS_XI39/MM4097_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2177 XI39/NET10638 N_NET264_XI39/MM2177_g N_VSS_XI39/MM2177_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4098 N_NET0380_XI39/MM4098_d N_NET265_XI39/MM4098_g N_VSS_XI39/MM4098_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2241 XI39/NET10390 N_NET396_XI39/MM2241_g N_VSS_XI39/MM2241_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4099 N_NET0380_XI39/MM4099_d N_NET267_XI39/MM4099_g N_VSS_XI39/MM4099_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2288 XI39/NET10210 N_NET268_XI39/MM2288_g N_VSS_XI39/MM2288_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4100 N_NET0380_XI39/MM4100_d N_NET269_XI39/MM4100_g N_VSS_XI39/MM4100_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2113 XI39/NET9874 N_NET270_XI39/MM2113_g N_VSS_XI39/MM2113_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4101 N_NET0380_XI39/MM4101_d N_NET401_XI39/MM4101_g N_VSS_XI39/MM4101_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2160 XI39/NET9694 N_NET272_XI39/MM2160_g N_VSS_XI39/MM2160_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4102 N_NET0380_XI39/MM4102_d N_NET273_XI39/MM4102_g N_VSS_XI39/MM4102_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2096 XI39/NET9946 N_NET404_XI39/MM2096_g N_VSS_XI39/MM2096_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4096 N_NET0380_XI39/MM4096_d N_NET405_XI39/MM4096_g N_VSS_XI39/MM4096_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM14 XI39/NET10098 N_NET0390_XI39/MM14_g N_VSS_XI39/MM14_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI29/XI0/MM39 N_NET0380_XI29/XI0/MM39_d N_XI29/XI0/NET195_XI29/XI0/MM39_g
+ N_NET064_XI29/XI0/MM39_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI29/XI0/XI8/MM1 N_XI29/XI0/NET195_XI29/XI0/XI8/MM1_d
+ N_NET470_XI29/XI0/XI8/MM1_g N_VSS_XI29/XI0/XI8/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI29/XI0/MM40 N_NET474_XI29/XI0/MM40_d N_XI29/XI0/NET199_XI29/XI0/MM40_g
+ N_NET064_XI29/XI0/MM40_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI29/XI0/XI9/MM1 N_XI29/XI0/NET199_XI29/XI0/XI9/MM1_d
+ N_NET469_XI29/XI0/XI9/MM1_g N_VSS_XI29/XI0/XI9/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI39/MM3408 XI39/NET5590 N_NET0133_XI39/MM3408_g N_VSS_XI39/MM3408_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3406 N_NET474_XI39/MM3406_d N_NET280_XI39/MM3406_g N_VSS_XI39/MM3406_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3423 XI39/NET5530 N_NET281_XI39/MM3423_g N_VSS_XI39/MM3423_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3440 N_NET474_XI39/MM3440_d N_NET282_XI39/MM3440_g N_VSS_XI39/MM3440_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3360 XI39/NET5782 N_NET153_XI39/MM3360_g N_VSS_XI39/MM3360_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3377 N_NET474_XI39/MM3377_d N_NET284_XI39/MM3377_g N_VSS_XI39/MM3377_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3345 XI39/NET3542 N_NET285_XI39/MM3345_g N_VSS_XI39/MM3345_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3342 N_NET474_XI39/MM3342_d N_NET286_XI39/MM3342_g N_VSS_XI39/MM3342_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3487 XI39/NET5274 N_NET287_XI39/MM3487_g N_VSS_XI39/MM3487_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3504 N_NET474_XI39/MM3504_d N_NET158_XI39/MM3504_g N_VSS_XI39/MM3504_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3472 XI39/NET5334 N_NET159_XI39/MM3472_g N_VSS_XI39/MM3472_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3469 N_NET474_XI39/MM3469_d N_NET160_XI39/MM3469_g N_VSS_XI39/MM3469_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3536 XI39/NET5078 N_NET291_XI39/MM3536_g N_VSS_XI39/MM3536_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3533 N_NET474_XI39/MM3533_d N_NET162_XI39/MM3533_g N_VSS_XI39/MM3533_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3551 XI39/NET5018 N_NET293_XI39/MM3551_g N_VSS_XI39/MM3551_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3568 N_NET474_XI39/MM3568_d N_NET294_XI39/MM3568_g N_VSS_XI39/MM3568_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3232 XI39/NET3994 N_NET295_XI39/MM3232_g N_VSS_XI39/MM3232_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3249 N_NET474_XI39/MM3249_d N_NET296_XI39/MM3249_g N_VSS_XI39/MM3249_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3217 XI39/NET4054 N_NET297_XI39/MM3217_g N_VSS_XI39/MM3217_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3214 N_NET474_XI39/MM3214_d N_NET298_XI39/MM3214_g N_VSS_XI39/MM3214_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3281 XI39/NET3798 N_NET299_XI39/MM3281_g N_VSS_XI39/MM3281_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3278 N_NET474_XI39/MM3278_d N_NET170_XI39/MM3278_g N_VSS_XI39/MM3278_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3296 XI39/NET3738 N_NET171_XI39/MM3296_g N_VSS_XI39/MM3296_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3313 N_NET474_XI39/MM3313_d N_NET172_XI39/MM3313_g N_VSS_XI39/MM3313_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3153 XI39/NET4310 N_NET303_XI39/MM3153_g N_VSS_XI39/MM3153_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3150 N_NET474_XI39/MM3150_d N_NET304_XI39/MM3150_g N_VSS_XI39/MM3150_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3168 XI39/NET4250 N_NET305_XI39/MM3168_g N_VSS_XI39/MM3168_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3185 N_NET474_XI39/MM3185_d N_NET306_XI39/MM3185_g N_VSS_XI39/MM3185_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3104 XI39/NET4506 N_NET307_XI39/MM3104_g N_VSS_XI39/MM3104_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3121 N_NET474_XI39/MM3121_d N_NET308_XI39/MM3121_g N_VSS_XI39/MM3121_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3089 XI39/NET4566 N_NET309_XI39/MM3089_g N_VSS_XI39/MM3089_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3086 N_NET474_XI39/MM3086_d N_NET310_XI39/MM3086_g N_VSS_XI39/MM3086_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3995 XI39/NET7338 N_NET311_XI39/MM3995_g N_VSS_XI39/MM3995_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3850 N_NET474_XI39/MM3850_d N_NET312_XI39/MM3850_g N_VSS_XI39/MM3850_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3980 XI39/NET7398 N_NET313_XI39/MM3980_g N_VSS_XI39/MM3980_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3977 N_NET474_XI39/MM3977_d N_NET314_XI39/MM3977_g N_VSS_XI39/MM3977_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3882 XI39/NET5994 N_NET315_XI39/MM3882_g N_VSS_XI39/MM3882_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3879 N_NET474_XI39/MM3879_d N_NET316_XI39/MM3879_g N_VSS_XI39/MM3879_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3897 XI39/NET5934 N_NET317_XI39/MM3897_g N_VSS_XI39/MM3897_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3914 N_NET474_XI39/MM3914_d N_NET318_XI39/MM3914_g N_VSS_XI39/MM3914_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4060 XI39/NET7078 N_NET319_XI39/MM4060_g N_VSS_XI39/MM4060_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4057 N_NET474_XI39/MM4057_d N_NET320_XI39/MM4057_g N_VSS_XI39/MM4057_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3935 XI39/NET7578 N_NET321_XI39/MM3935_g N_VSS_XI39/MM3935_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3948 N_NET474_XI39/MM3948_d N_NET192_XI39/MM3948_g N_VSS_XI39/MM3948_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4011 XI39/NET7274 N_NET193_XI39/MM4011_g N_VSS_XI39/MM4011_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4028 N_NET474_XI39/MM4028_d N_NET194_XI39/MM4028_g N_VSS_XI39/MM4028_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4002 XI39/NET7310 N_NET195_XI39/MM4002_g N_VSS_XI39/MM4002_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4087 N_NET474_XI39/MM4087_d N_NET196_XI39/MM4087_g N_VSS_XI39/MM4087_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3792 XI39/NET6354 N_NET197_XI39/MM3792_g N_VSS_XI39/MM3792_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3789 N_NET474_XI39/MM3789_d N_NET198_XI39/MM3789_g N_VSS_XI39/MM3789_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3807 XI39/NET6294 N_NET199_XI39/MM3807_g N_VSS_XI39/MM3807_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3824 N_NET474_XI39/MM3824_d N_NET200_XI39/MM3824_g N_VSS_XI39/MM3824_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3743 XI39/NET6550 N_NET331_XI39/MM3743_g N_VSS_XI39/MM3743_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3760 N_NET474_XI39/MM3760_d N_NET332_XI39/MM3760_g N_VSS_XI39/MM3760_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3728 XI39/NET6610 N_NET203_XI39/MM3728_g N_VSS_XI39/MM3728_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3725 N_NET474_XI39/MM3725_d N_NET204_XI39/MM3725_g N_VSS_XI39/MM3725_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3615 XI39/NET4762 N_NET205_XI39/MM3615_g N_VSS_XI39/MM3615_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3632 N_NET474_XI39/MM3632_d N_NET206_XI39/MM3632_g N_VSS_XI39/MM3632_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3600 XI39/NET4822 N_NET207_XI39/MM3600_g N_VSS_XI39/MM3600_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3597 N_NET474_XI39/MM3597_d N_NET338_XI39/MM3597_g N_VSS_XI39/MM3597_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3664 XI39/NET6866 N_NET339_XI39/MM3664_g N_VSS_XI39/MM3664_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3661 N_NET474_XI39/MM3661_d N_NET340_XI39/MM3661_g N_VSS_XI39/MM3661_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3680 XI39/NET6802 N_NET211_XI39/MM3680_g N_VSS_XI39/MM3680_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3689 N_NET474_XI39/MM3689_d N_NET212_XI39/MM3689_g N_VSS_XI39/MM3689_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2720 XI39/NET8982 N_NET214_XI39/MM2720_g N_VSS_XI39/MM2720_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2737 N_NET474_XI39/MM2737_d N_NET215_XI39/MM2737_g N_VSS_XI39/MM2737_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2705 XI39/NET9042 N_NET216_XI39/MM2705_g N_VSS_XI39/MM2705_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2702 N_NET474_XI39/MM2702_d N_NET346_XI39/MM2702_g N_VSS_XI39/MM2702_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2769 XI39/NET8790 N_NET347_XI39/MM2769_g N_VSS_XI39/MM2769_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2766 N_NET474_XI39/MM2766_d N_NET348_XI39/MM2766_g N_VSS_XI39/MM2766_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2784 XI39/NET8730 N_NET349_XI39/MM2784_g N_VSS_XI39/MM2784_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2801 N_NET474_XI39/MM2801_d N_NET350_XI39/MM2801_g N_VSS_XI39/MM2801_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2641 XI39/NET9298 N_NET351_XI39/MM2641_g N_VSS_XI39/MM2641_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2638 N_NET474_XI39/MM2638_d N_NET352_XI39/MM2638_g N_VSS_XI39/MM2638_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2656 XI39/NET9238 N_NET224_XI39/MM2656_g N_VSS_XI39/MM2656_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2673 N_NET474_XI39/MM2673_d N_NET225_XI39/MM2673_g N_VSS_XI39/MM2673_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2592 XI39/NET9494 N_NET226_XI39/MM2592_g N_VSS_XI39/MM2592_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2609 N_NET474_XI39/MM2609_d N_NET356_XI39/MM2609_g N_VSS_XI39/MM2609_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2577 XI39/NET9554 N_NET357_XI39/MM2577_g N_VSS_XI39/MM2577_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2574 N_NET474_XI39/MM2574_d N_NET358_XI39/MM2574_g N_VSS_XI39/MM2574_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2897 XI39/NET8278 N_NET230_XI39/MM2897_g N_VSS_XI39/MM2897_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2894 N_NET474_XI39/MM2894_d N_NET360_XI39/MM2894_g N_VSS_XI39/MM2894_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2912 XI39/NET8218 N_NET361_XI39/MM2912_g N_VSS_XI39/MM2912_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2929 N_NET474_XI39/MM2929_d N_NET233_XI39/MM2929_g N_VSS_XI39/MM2929_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2848 XI39/NET8474 N_NET234_XI39/MM2848_g N_VSS_XI39/MM2848_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2865 N_NET474_XI39/MM2865_d N_NET235_XI39/MM2865_g N_VSS_XI39/MM2865_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2833 XI39/NET8534 N_NET365_XI39/MM2833_g N_VSS_XI39/MM2833_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2830 N_NET474_XI39/MM2830_d N_NET366_XI39/MM2830_g N_VSS_XI39/MM2830_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2976 XI39/NET7962 N_NET367_XI39/MM2976_g N_VSS_XI39/MM2976_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2993 N_NET474_XI39/MM2993_d N_NET368_XI39/MM2993_g N_VSS_XI39/MM2993_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2961 XI39/NET8022 N_NET369_XI39/MM2961_g N_VSS_XI39/MM2961_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2958 N_NET474_XI39/MM2958_d N_NET370_XI39/MM2958_g N_VSS_XI39/MM2958_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3025 XI39/NET7766 N_NET371_XI39/MM3025_g N_VSS_XI39/MM3025_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3022 N_NET474_XI39/MM3022_d N_NET242_XI39/MM3022_g N_VSS_XI39/MM3022_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3040 XI39/NET7706 N_NET373_XI39/MM3040_g N_VSS_XI39/MM3040_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3057 N_NET474_XI39/MM3057_d N_NET244_XI39/MM3057_g N_VSS_XI39/MM3057_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2395 XI39/NET11290 N_NET375_XI39/MM2395_g N_VSS_XI39/MM2395_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2382 N_NET474_XI39/MM2382_d N_NET376_XI39/MM2382_g N_VSS_XI39/MM2382_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2400 XI39/NET11270 N_NET377_XI39/MM2400_g N_VSS_XI39/MM2400_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2417 N_NET474_XI39/MM2417_d N_NET378_XI39/MM2417_g N_VSS_XI39/MM2417_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2336 XI39/NET10878 N_NET379_XI39/MM2336_g N_VSS_XI39/MM2336_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2353 N_NET474_XI39/MM2353_d N_NET380_XI39/MM2353_g N_VSS_XI39/MM2353_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2321 XI39/NET10938 N_NET381_XI39/MM2321_g N_VSS_XI39/MM2321_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2318 N_NET474_XI39/MM2318_d N_NET382_XI39/MM2318_g N_VSS_XI39/MM2318_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2466 XI39/NET11582 N_NET383_XI39/MM2466_g N_VSS_XI39/MM2466_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2481 N_NET474_XI39/MM2481_d N_NET384_XI39/MM2481_g N_VSS_XI39/MM2481_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2449 XI39/NET11074 N_NET385_XI39/MM2449_g N_VSS_XI39/MM2449_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2446 N_NET474_XI39/MM2446_d N_NET256_XI39/MM2446_g N_VSS_XI39/MM2446_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2513 XI39/NET11394 N_NET387_XI39/MM2513_g N_VSS_XI39/MM2513_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2510 N_NET474_XI39/MM2510_d N_NET388_XI39/MM2510_g N_VSS_XI39/MM2510_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2538 XI39/NET11670 N_NET389_XI39/MM2538_g N_VSS_XI39/MM2538_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2545 N_NET474_XI39/MM2545_d N_NET390_XI39/MM2545_g N_VSS_XI39/MM2545_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2208 XI39/NET10518 N_NET391_XI39/MM2208_g N_VSS_XI39/MM2208_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2225 N_NET474_XI39/MM2225_d N_NET262_XI39/MM2225_g N_VSS_XI39/MM2225_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2193 XI39/NET10578 N_NET263_XI39/MM2193_g N_VSS_XI39/MM2193_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2190 N_NET474_XI39/MM2190_d N_NET264_XI39/MM2190_g N_VSS_XI39/MM2190_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2257 XI39/NET10330 N_NET265_XI39/MM2257_g N_VSS_XI39/MM2257_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2254 N_NET474_XI39/MM2254_d N_NET396_XI39/MM2254_g N_VSS_XI39/MM2254_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2272 XI39/NET10270 N_NET267_XI39/MM2272_g N_VSS_XI39/MM2272_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2289 N_NET474_XI39/MM2289_d N_NET268_XI39/MM2289_g N_VSS_XI39/MM2289_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2129 XI39/NET9814 N_NET269_XI39/MM2129_g N_VSS_XI39/MM2129_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2126 N_NET474_XI39/MM2126_d N_NET270_XI39/MM2126_g N_VSS_XI39/MM2126_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2144 XI39/NET9754 N_NET401_XI39/MM2144_g N_VSS_XI39/MM2144_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2161 N_NET474_XI39/MM2161_d N_NET272_XI39/MM2161_g N_VSS_XI39/MM2161_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2080 XI39/NET10006 N_NET273_XI39/MM2080_g N_VSS_XI39/MM2080_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2097 N_NET474_XI39/MM2097_d N_NET404_XI39/MM2097_g N_VSS_XI39/MM2097_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2079 XI39/NET10130 N_NET405_XI39/MM2079_g N_VSS_XI39/MM2079_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM1 N_NET474_XI39/MM1_d N_NET0390_XI39/MM1_g N_VSS_XI39/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI57/XI1/MM7 N_XI57/XI1/NET1_XI57/XI1/MM7_d N_NET065_XI57/XI1/MM7_g
+ N_XI57/XI1/NET9_XI57/XI1/MM7_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=1.2e-06 AD=4.5e-13 AS=6e-13 PD=7.5e-07 PS=2.2e-06
mXI57/XI1/MM5 N_XI57/NET12_XI57/XI1/MM5_d N_NET061_XI57/XI1/MM5_g
+ N_XI57/XI1/NET1_XI57/XI1/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=1.2e-06 AD=6.06e-13 AS=4.5e-13 PD=2.21e-06 PS=7.5e-07
mXI57/XI1/MM4 N_NET061_XI57/XI1/MM4_d N_XI57/NET12_XI57/XI1/MM4_g
+ N_XI57/XI1/NET20_XI57/XI1/MM4_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18
+ L=1.8e-07 W=1.2e-06 AD=6.06e-13 AS=4.5e-13 PD=2.21e-06 PS=7.5e-07
mXI57/XI1/MM6 N_XI57/XI1/NET20_XI57/XI1/MM6_d N_VREF_XI57/XI1/MM6_g
+ N_XI57/XI1/NET9_XI57/XI1/MM6_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=1.2e-06 AD=4.5e-13 AS=6e-13 PD=7.5e-07 PS=2.2e-06
mXI57/XI1/MM8 N_XI57/XI1/NET9_XI57/XI1/MM8_d N_NET068_XI57/XI1/MM8_g
+ N_VSS_XI57/XI1/MM8_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI29/XI0/MM41 N_NET475_XI29/XI0/MM41_d N_XI29/XI0/NET223_XI29/XI0/MM41_g
+ N_NET064_XI29/XI0/MM41_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI29/XI0/XI10/MM1 N_XI29/XI0/NET223_XI29/XI0/XI10/MM1_d
+ N_NET468_XI29/XI0/XI10/MM1_g N_VSS_XI29/XI0/XI10/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI29/XI0/MM42 N_NET476_XI29/XI0/MM42_d N_XI29/XI0/NET215_XI29/XI0/MM42_g
+ N_NET064_XI29/XI0/MM42_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI29/XI0/XI11/MM1 N_XI29/XI0/NET215_XI29/XI0/XI11/MM1_d
+ N_NET467_XI29/XI0/XI11/MM1_g N_VSS_XI29/XI0/XI11/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI39/MM3409 N_NET475_XI39/MM3409_d N_NET0133_XI39/MM3409_g N_VSS_XI39/MM3409_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3407 XI39/NET5594 N_NET280_XI39/MM3407_g N_VSS_XI39/MM3407_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3436 N_NET475_XI39/MM3436_d N_NET281_XI39/MM3436_g N_VSS_XI39/MM3436_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3453 XI39/NET5410 N_NET282_XI39/MM3453_g N_VSS_XI39/MM3453_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3373 N_NET475_XI39/MM3373_d N_NET153_XI39/MM3373_g N_VSS_XI39/MM3373_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3390 XI39/NET5662 N_NET284_XI39/MM3390_g N_VSS_XI39/MM3390_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3346 N_NET475_XI39/MM3346_d N_NET285_XI39/MM3346_g N_VSS_XI39/MM3346_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3339 XI39/NET3566 N_NET286_XI39/MM3339_g N_VSS_XI39/MM3339_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3500 N_NET475_XI39/MM3500_d N_NET287_XI39/MM3500_g N_VSS_XI39/MM3500_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3517 XI39/NET5154 N_NET158_XI39/MM3517_g N_VSS_XI39/MM3517_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3473 N_NET475_XI39/MM3473_d N_NET159_XI39/MM3473_g N_VSS_XI39/MM3473_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3470 XI39/NET5342 N_NET160_XI39/MM3470_g N_VSS_XI39/MM3470_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3537 N_NET475_XI39/MM3537_d N_NET291_XI39/MM3537_g N_VSS_XI39/MM3537_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3534 XI39/NET5086 N_NET162_XI39/MM3534_g N_VSS_XI39/MM3534_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3564 N_NET475_XI39/MM3564_d N_NET293_XI39/MM3564_g N_VSS_XI39/MM3564_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3581 XI39/NET4898 N_NET294_XI39/MM3581_g N_VSS_XI39/MM3581_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3245 N_NET475_XI39/MM3245_d N_NET295_XI39/MM3245_g N_VSS_XI39/MM3245_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3262 XI39/NET3874 N_NET296_XI39/MM3262_g N_VSS_XI39/MM3262_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3218 N_NET475_XI39/MM3218_d N_NET297_XI39/MM3218_g N_VSS_XI39/MM3218_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3215 XI39/NET4062 N_NET298_XI39/MM3215_g N_VSS_XI39/MM3215_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3282 N_NET475_XI39/MM3282_d N_NET299_XI39/MM3282_g N_VSS_XI39/MM3282_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3279 XI39/NET3806 N_NET170_XI39/MM3279_g N_VSS_XI39/MM3279_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3309 N_NET475_XI39/MM3309_d N_NET171_XI39/MM3309_g N_VSS_XI39/MM3309_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3326 XI39/NET3618 N_NET172_XI39/MM3326_g N_VSS_XI39/MM3326_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3154 N_NET475_XI39/MM3154_d N_NET303_XI39/MM3154_g N_VSS_XI39/MM3154_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3151 XI39/NET4318 N_NET304_XI39/MM3151_g N_VSS_XI39/MM3151_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3181 N_NET475_XI39/MM3181_d N_NET305_XI39/MM3181_g N_VSS_XI39/MM3181_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3198 XI39/NET4130 N_NET306_XI39/MM3198_g N_VSS_XI39/MM3198_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3117 N_NET475_XI39/MM3117_d N_NET307_XI39/MM3117_g N_VSS_XI39/MM3117_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3134 XI39/NET4386 N_NET308_XI39/MM3134_g N_VSS_XI39/MM3134_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3090 N_NET475_XI39/MM3090_d N_NET309_XI39/MM3090_g N_VSS_XI39/MM3090_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3087 XI39/NET4574 N_NET310_XI39/MM3087_g N_VSS_XI39/MM3087_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3846 N_NET475_XI39/MM3846_d N_NET311_XI39/MM3846_g N_VSS_XI39/MM3846_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3863 XI39/NET6070 N_NET312_XI39/MM3863_g N_VSS_XI39/MM3863_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3981 N_NET475_XI39/MM3981_d N_NET313_XI39/MM3981_g N_VSS_XI39/MM3981_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3978 XI39/NET7406 N_NET314_XI39/MM3978_g N_VSS_XI39/MM3978_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3883 N_NET475_XI39/MM3883_d N_NET315_XI39/MM3883_g N_VSS_XI39/MM3883_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3880 XI39/NET6002 N_NET316_XI39/MM3880_g N_VSS_XI39/MM3880_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3910 N_NET475_XI39/MM3910_d N_NET317_XI39/MM3910_g N_VSS_XI39/MM3910_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3927 XI39/NET5814 N_NET318_XI39/MM3927_g N_VSS_XI39/MM3927_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4061 N_NET475_XI39/MM4061_d N_NET319_XI39/MM4061_g N_VSS_XI39/MM4061_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4058 XI39/NET7086 N_NET320_XI39/MM4058_g N_VSS_XI39/MM4058_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3944 N_NET475_XI39/MM3944_d N_NET321_XI39/MM3944_g N_VSS_XI39/MM3944_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3961 XI39/NET7474 N_NET192_XI39/MM3961_g N_VSS_XI39/MM3961_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4024 N_NET475_XI39/MM4024_d N_NET193_XI39/MM4024_g N_VSS_XI39/MM4024_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4041 XI39/NET7154 N_NET194_XI39/MM4041_g N_VSS_XI39/MM4041_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4091 N_NET475_XI39/MM4091_d N_NET195_XI39/MM4091_g N_VSS_XI39/MM4091_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4088 XI39/NET6966 N_NET196_XI39/MM4088_g N_VSS_XI39/MM4088_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3793 N_NET475_XI39/MM3793_d N_NET197_XI39/MM3793_g N_VSS_XI39/MM3793_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3790 XI39/NET6362 N_NET198_XI39/MM3790_g N_VSS_XI39/MM3790_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3820 N_NET475_XI39/MM3820_d N_NET199_XI39/MM3820_g N_VSS_XI39/MM3820_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3837 XI39/NET6174 N_NET200_XI39/MM3837_g N_VSS_XI39/MM3837_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3756 N_NET475_XI39/MM3756_d N_NET331_XI39/MM3756_g N_VSS_XI39/MM3756_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3773 XI39/NET6430 N_NET332_XI39/MM3773_g N_VSS_XI39/MM3773_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3729 N_NET475_XI39/MM3729_d N_NET203_XI39/MM3729_g N_VSS_XI39/MM3729_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3726 XI39/NET6618 N_NET204_XI39/MM3726_g N_VSS_XI39/MM3726_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3628 N_NET475_XI39/MM3628_d N_NET205_XI39/MM3628_g N_VSS_XI39/MM3628_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3645 XI39/NET4642 N_NET206_XI39/MM3645_g N_VSS_XI39/MM3645_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3601 N_NET475_XI39/MM3601_d N_NET207_XI39/MM3601_g N_VSS_XI39/MM3601_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3598 XI39/NET4830 N_NET338_XI39/MM3598_g N_VSS_XI39/MM3598_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3665 N_NET475_XI39/MM3665_d N_NET339_XI39/MM3665_g N_VSS_XI39/MM3665_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3662 XI39/NET6874 N_NET340_XI39/MM3662_g N_VSS_XI39/MM3662_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3681 N_NET475_XI39/MM3681_d N_NET211_XI39/MM3681_g N_VSS_XI39/MM3681_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3702 XI39/NET6714 N_NET212_XI39/MM3702_g N_VSS_XI39/MM3702_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2733 N_NET475_XI39/MM2733_d N_NET214_XI39/MM2733_g N_VSS_XI39/MM2733_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2750 XI39/NET8866 N_NET215_XI39/MM2750_g N_VSS_XI39/MM2750_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2706 N_NET475_XI39/MM2706_d N_NET216_XI39/MM2706_g N_VSS_XI39/MM2706_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2703 XI39/NET9050 N_NET346_XI39/MM2703_g N_VSS_XI39/MM2703_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2770 N_NET475_XI39/MM2770_d N_NET347_XI39/MM2770_g N_VSS_XI39/MM2770_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2767 XI39/NET8798 N_NET348_XI39/MM2767_g N_VSS_XI39/MM2767_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2797 N_NET475_XI39/MM2797_d N_NET349_XI39/MM2797_g N_VSS_XI39/MM2797_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2814 XI39/NET8610 N_NET350_XI39/MM2814_g N_VSS_XI39/MM2814_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2642 N_NET475_XI39/MM2642_d N_NET351_XI39/MM2642_g N_VSS_XI39/MM2642_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2639 XI39/NET9306 N_NET352_XI39/MM2639_g N_VSS_XI39/MM2639_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2669 N_NET475_XI39/MM2669_d N_NET224_XI39/MM2669_g N_VSS_XI39/MM2669_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2686 XI39/NET9118 N_NET225_XI39/MM2686_g N_VSS_XI39/MM2686_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2605 N_NET475_XI39/MM2605_d N_NET226_XI39/MM2605_g N_VSS_XI39/MM2605_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2622 XI39/NET9374 N_NET356_XI39/MM2622_g N_VSS_XI39/MM2622_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2578 N_NET475_XI39/MM2578_d N_NET357_XI39/MM2578_g N_VSS_XI39/MM2578_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2575 XI39/NET9562 N_NET358_XI39/MM2575_g N_VSS_XI39/MM2575_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2898 N_NET475_XI39/MM2898_d N_NET230_XI39/MM2898_g N_VSS_XI39/MM2898_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2895 XI39/NET8286 N_NET360_XI39/MM2895_g N_VSS_XI39/MM2895_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2925 N_NET475_XI39/MM2925_d N_NET361_XI39/MM2925_g N_VSS_XI39/MM2925_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2942 XI39/NET8098 N_NET233_XI39/MM2942_g N_VSS_XI39/MM2942_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2861 N_NET475_XI39/MM2861_d N_NET234_XI39/MM2861_g N_VSS_XI39/MM2861_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2878 XI39/NET8354 N_NET235_XI39/MM2878_g N_VSS_XI39/MM2878_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2834 N_NET475_XI39/MM2834_d N_NET365_XI39/MM2834_g N_VSS_XI39/MM2834_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2831 XI39/NET8542 N_NET366_XI39/MM2831_g N_VSS_XI39/MM2831_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2989 N_NET475_XI39/MM2989_d N_NET367_XI39/MM2989_g N_VSS_XI39/MM2989_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3006 XI39/NET7842 N_NET368_XI39/MM3006_g N_VSS_XI39/MM3006_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2962 N_NET475_XI39/MM2962_d N_NET369_XI39/MM2962_g N_VSS_XI39/MM2962_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2959 XI39/NET8030 N_NET370_XI39/MM2959_g N_VSS_XI39/MM2959_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3026 N_NET475_XI39/MM3026_d N_NET371_XI39/MM3026_g N_VSS_XI39/MM3026_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3023 XI39/NET7774 N_NET242_XI39/MM3023_g N_VSS_XI39/MM3023_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3053 N_NET475_XI39/MM3053_d N_NET373_XI39/MM3053_g N_VSS_XI39/MM3053_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3070 XI39/NET7586 N_NET244_XI39/MM3070_g N_VSS_XI39/MM3070_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2386 N_NET475_XI39/MM2386_d N_NET375_XI39/MM2386_g N_VSS_XI39/MM2386_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2383 XI39/NET10690 N_NET376_XI39/MM2383_g N_VSS_XI39/MM2383_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2413 N_NET475_XI39/MM2413_d N_NET377_XI39/MM2413_g N_VSS_XI39/MM2413_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2430 XI39/NET11150 N_NET378_XI39/MM2430_g N_VSS_XI39/MM2430_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2349 N_NET475_XI39/MM2349_d N_NET379_XI39/MM2349_g N_VSS_XI39/MM2349_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2366 XI39/NET10758 N_NET380_XI39/MM2366_g N_VSS_XI39/MM2366_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2322 N_NET475_XI39/MM2322_d N_NET381_XI39/MM2322_g N_VSS_XI39/MM2322_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2319 XI39/NET10946 N_NET382_XI39/MM2319_g N_VSS_XI39/MM2319_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2477 N_NET475_XI39/MM2477_d N_NET383_XI39/MM2477_g N_VSS_XI39/MM2477_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2494 XI39/NET11470 N_NET384_XI39/MM2494_g N_VSS_XI39/MM2494_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2450 N_NET475_XI39/MM2450_d N_NET385_XI39/MM2450_g N_VSS_XI39/MM2450_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2447 XI39/NET11082 N_NET256_XI39/MM2447_g N_VSS_XI39/MM2447_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2514 N_NET475_XI39/MM2514_d N_NET387_XI39/MM2514_g N_VSS_XI39/MM2514_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2511 XI39/NET11402 N_NET388_XI39/MM2511_g N_VSS_XI39/MM2511_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2541 N_NET475_XI39/MM2541_d N_NET389_XI39/MM2541_g N_VSS_XI39/MM2541_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2558 XI39/NET11590 N_NET390_XI39/MM2558_g N_VSS_XI39/MM2558_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2221 N_NET475_XI39/MM2221_d N_NET391_XI39/MM2221_g N_VSS_XI39/MM2221_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2238 XI39/NET10402 N_NET262_XI39/MM2238_g N_VSS_XI39/MM2238_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2194 N_NET475_XI39/MM2194_d N_NET263_XI39/MM2194_g N_VSS_XI39/MM2194_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2191 XI39/NET10582 N_NET264_XI39/MM2191_g N_VSS_XI39/MM2191_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2258 N_NET475_XI39/MM2258_d N_NET265_XI39/MM2258_g N_VSS_XI39/MM2258_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2255 XI39/NET10334 N_NET396_XI39/MM2255_g N_VSS_XI39/MM2255_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2285 N_NET475_XI39/MM2285_d N_NET267_XI39/MM2285_g N_VSS_XI39/MM2285_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2302 XI39/NET10154 N_NET268_XI39/MM2302_g N_VSS_XI39/MM2302_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2130 N_NET475_XI39/MM2130_d N_NET269_XI39/MM2130_g N_VSS_XI39/MM2130_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2127 XI39/NET9818 N_NET270_XI39/MM2127_g N_VSS_XI39/MM2127_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2157 N_NET475_XI39/MM2157_d N_NET401_XI39/MM2157_g N_VSS_XI39/MM2157_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2174 XI39/NET9638 N_NET272_XI39/MM2174_g N_VSS_XI39/MM2174_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2093 N_NET475_XI39/MM2093_d N_NET273_XI39/MM2093_g N_VSS_XI39/MM2093_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2110 XI39/NET9890 N_NET404_XI39/MM2110_g N_VSS_XI39/MM2110_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2066 N_NET475_XI39/MM2066_d N_NET405_XI39/MM2066_g N_VSS_XI39/MM2066_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM6 XI39/NET10066 N_NET0390_XI39/MM6_g N_VSS_XI39/MM6_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3416 XI39/NET5558 N_NET0133_XI39/MM3416_g N_VSS_XI39/MM3416_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3404 N_NET476_XI39/MM3404_d N_NET280_XI39/MM3404_g N_VSS_XI39/MM3404_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3435 XI39/NET5482 N_NET281_XI39/MM3435_g N_VSS_XI39/MM3435_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3442 N_NET476_XI39/MM3442_d N_NET282_XI39/MM3442_g N_VSS_XI39/MM3442_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3372 XI39/NET5734 N_NET153_XI39/MM3372_g N_VSS_XI39/MM3372_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3379 N_NET476_XI39/MM3379_d N_NET284_XI39/MM3379_g N_VSS_XI39/MM3379_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3357 XI39/NET3494 N_NET285_XI39/MM3357_g N_VSS_XI39/MM3357_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3340 N_NET476_XI39/MM3340_d N_NET286_XI39/MM3340_g N_VSS_XI39/MM3340_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3499 XI39/NET5226 N_NET287_XI39/MM3499_g N_VSS_XI39/MM3499_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3506 N_NET476_XI39/MM3506_d N_NET158_XI39/MM3506_g N_VSS_XI39/MM3506_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3484 XI39/NET5286 N_NET159_XI39/MM3484_g N_VSS_XI39/MM3484_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3467 N_NET476_XI39/MM3467_d N_NET160_XI39/MM3467_g N_VSS_XI39/MM3467_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3548 XI39/NET5030 N_NET291_XI39/MM3548_g N_VSS_XI39/MM3548_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3531 N_NET476_XI39/MM3531_d N_NET162_XI39/MM3531_g N_VSS_XI39/MM3531_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3563 XI39/NET4970 N_NET293_XI39/MM3563_g N_VSS_XI39/MM3563_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3570 N_NET476_XI39/MM3570_d N_NET294_XI39/MM3570_g N_VSS_XI39/MM3570_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3244 XI39/NET3946 N_NET295_XI39/MM3244_g N_VSS_XI39/MM3244_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3251 N_NET476_XI39/MM3251_d N_NET296_XI39/MM3251_g N_VSS_XI39/MM3251_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3229 XI39/NET4006 N_NET297_XI39/MM3229_g N_VSS_XI39/MM3229_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3212 N_NET476_XI39/MM3212_d N_NET298_XI39/MM3212_g N_VSS_XI39/MM3212_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3293 XI39/NET3750 N_NET299_XI39/MM3293_g N_VSS_XI39/MM3293_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3276 N_NET476_XI39/MM3276_d N_NET170_XI39/MM3276_g N_VSS_XI39/MM3276_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3308 XI39/NET3690 N_NET171_XI39/MM3308_g N_VSS_XI39/MM3308_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3315 N_NET476_XI39/MM3315_d N_NET172_XI39/MM3315_g N_VSS_XI39/MM3315_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3165 XI39/NET4262 N_NET303_XI39/MM3165_g N_VSS_XI39/MM3165_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3148 N_NET476_XI39/MM3148_d N_NET304_XI39/MM3148_g N_VSS_XI39/MM3148_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3180 XI39/NET4202 N_NET305_XI39/MM3180_g N_VSS_XI39/MM3180_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3187 N_NET476_XI39/MM3187_d N_NET306_XI39/MM3187_g N_VSS_XI39/MM3187_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3116 XI39/NET4458 N_NET307_XI39/MM3116_g N_VSS_XI39/MM3116_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3123 N_NET476_XI39/MM3123_d N_NET308_XI39/MM3123_g N_VSS_XI39/MM3123_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3101 XI39/NET4518 N_NET309_XI39/MM3101_g N_VSS_XI39/MM3101_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3084 N_NET476_XI39/MM3084_d N_NET310_XI39/MM3084_g N_VSS_XI39/MM3084_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3845 XI39/NET6142 N_NET311_XI39/MM3845_g N_VSS_XI39/MM3845_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3852 N_NET476_XI39/MM3852_d N_NET312_XI39/MM3852_g N_VSS_XI39/MM3852_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3992 XI39/NET7350 N_NET313_XI39/MM3992_g N_VSS_XI39/MM3992_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3975 N_NET476_XI39/MM3975_d N_NET314_XI39/MM3975_g N_VSS_XI39/MM3975_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3894 XI39/NET5946 N_NET315_XI39/MM3894_g N_VSS_XI39/MM3894_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3877 N_NET476_XI39/MM3877_d N_NET316_XI39/MM3877_g N_VSS_XI39/MM3877_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3909 XI39/NET5886 N_NET317_XI39/MM3909_g N_VSS_XI39/MM3909_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3916 N_NET476_XI39/MM3916_d N_NET318_XI39/MM3916_g N_VSS_XI39/MM3916_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4072 XI39/NET7030 N_NET319_XI39/MM4072_g N_VSS_XI39/MM4072_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4055 N_NET476_XI39/MM4055_d N_NET320_XI39/MM4055_g N_VSS_XI39/MM4055_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3931 XI39/NET5798 N_NET321_XI39/MM3931_g N_VSS_XI39/MM3931_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3950 N_NET476_XI39/MM3950_d N_NET192_XI39/MM3950_g N_VSS_XI39/MM3950_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4023 XI39/NET7226 N_NET193_XI39/MM4023_g N_VSS_XI39/MM4023_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4030 N_NET476_XI39/MM4030_d N_NET194_XI39/MM4030_g N_VSS_XI39/MM4030_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4092 XI39/NET6950 N_NET195_XI39/MM4092_g N_VSS_XI39/MM4092_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4085 N_NET476_XI39/MM4085_d N_NET196_XI39/MM4085_g N_VSS_XI39/MM4085_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3804 XI39/NET6306 N_NET197_XI39/MM3804_g N_VSS_XI39/MM3804_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3787 N_NET476_XI39/MM3787_d N_NET198_XI39/MM3787_g N_VSS_XI39/MM3787_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3819 XI39/NET6246 N_NET199_XI39/MM3819_g N_VSS_XI39/MM3819_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3826 N_NET476_XI39/MM3826_d N_NET200_XI39/MM3826_g N_VSS_XI39/MM3826_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3755 XI39/NET6502 N_NET331_XI39/MM3755_g N_VSS_XI39/MM3755_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3762 N_NET476_XI39/MM3762_d N_NET332_XI39/MM3762_g N_VSS_XI39/MM3762_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3740 XI39/NET6562 N_NET203_XI39/MM3740_g N_VSS_XI39/MM3740_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3723 N_NET476_XI39/MM3723_d N_NET204_XI39/MM3723_g N_VSS_XI39/MM3723_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3627 XI39/NET4714 N_NET205_XI39/MM3627_g N_VSS_XI39/MM3627_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3634 N_NET476_XI39/MM3634_d N_NET206_XI39/MM3634_g N_VSS_XI39/MM3634_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3612 XI39/NET4774 N_NET207_XI39/MM3612_g N_VSS_XI39/MM3612_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3595 N_NET476_XI39/MM3595_d N_NET338_XI39/MM3595_g N_VSS_XI39/MM3595_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3676 XI39/NET6818 N_NET339_XI39/MM3676_g N_VSS_XI39/MM3676_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3659 N_NET476_XI39/MM3659_d N_NET340_XI39/MM3659_g N_VSS_XI39/MM3659_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3708 XI39/NET6690 N_NET211_XI39/MM3708_g N_VSS_XI39/MM3708_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3691 N_NET476_XI39/MM3691_d N_NET212_XI39/MM3691_g N_VSS_XI39/MM3691_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2732 XI39/NET8934 N_NET214_XI39/MM2732_g N_VSS_XI39/MM2732_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2739 N_NET476_XI39/MM2739_d N_NET215_XI39/MM2739_g N_VSS_XI39/MM2739_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2717 XI39/NET8994 N_NET216_XI39/MM2717_g N_VSS_XI39/MM2717_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2700 N_NET476_XI39/MM2700_d N_NET346_XI39/MM2700_g N_VSS_XI39/MM2700_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2781 XI39/NET8742 N_NET347_XI39/MM2781_g N_VSS_XI39/MM2781_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2764 N_NET476_XI39/MM2764_d N_NET348_XI39/MM2764_g N_VSS_XI39/MM2764_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2796 XI39/NET8682 N_NET349_XI39/MM2796_g N_VSS_XI39/MM2796_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2803 N_NET476_XI39/MM2803_d N_NET350_XI39/MM2803_g N_VSS_XI39/MM2803_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2653 XI39/NET9250 N_NET351_XI39/MM2653_g N_VSS_XI39/MM2653_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2636 N_NET476_XI39/MM2636_d N_NET352_XI39/MM2636_g N_VSS_XI39/MM2636_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2668 XI39/NET9190 N_NET224_XI39/MM2668_g N_VSS_XI39/MM2668_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2675 N_NET476_XI39/MM2675_d N_NET225_XI39/MM2675_g N_VSS_XI39/MM2675_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2604 XI39/NET9446 N_NET226_XI39/MM2604_g N_VSS_XI39/MM2604_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2611 N_NET476_XI39/MM2611_d N_NET356_XI39/MM2611_g N_VSS_XI39/MM2611_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2589 XI39/NET9506 N_NET357_XI39/MM2589_g N_VSS_XI39/MM2589_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2572 N_NET476_XI39/MM2572_d N_NET358_XI39/MM2572_g N_VSS_XI39/MM2572_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2909 XI39/NET8230 N_NET230_XI39/MM2909_g N_VSS_XI39/MM2909_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2892 N_NET476_XI39/MM2892_d N_NET360_XI39/MM2892_g N_VSS_XI39/MM2892_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2924 XI39/NET8170 N_NET361_XI39/MM2924_g N_VSS_XI39/MM2924_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2931 N_NET476_XI39/MM2931_d N_NET233_XI39/MM2931_g N_VSS_XI39/MM2931_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2860 XI39/NET8426 N_NET234_XI39/MM2860_g N_VSS_XI39/MM2860_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2867 N_NET476_XI39/MM2867_d N_NET235_XI39/MM2867_g N_VSS_XI39/MM2867_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2845 XI39/NET8486 N_NET365_XI39/MM2845_g N_VSS_XI39/MM2845_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2828 N_NET476_XI39/MM2828_d N_NET366_XI39/MM2828_g N_VSS_XI39/MM2828_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2988 XI39/NET7914 N_NET367_XI39/MM2988_g N_VSS_XI39/MM2988_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2995 N_NET476_XI39/MM2995_d N_NET368_XI39/MM2995_g N_VSS_XI39/MM2995_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2973 XI39/NET7974 N_NET369_XI39/MM2973_g N_VSS_XI39/MM2973_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2956 N_NET476_XI39/MM2956_d N_NET370_XI39/MM2956_g N_VSS_XI39/MM2956_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3037 XI39/NET7718 N_NET371_XI39/MM3037_g N_VSS_XI39/MM3037_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3020 N_NET476_XI39/MM3020_d N_NET242_XI39/MM3020_g N_VSS_XI39/MM3020_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3052 XI39/NET7658 N_NET373_XI39/MM3052_g N_VSS_XI39/MM3052_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3059 N_NET476_XI39/MM3059_d N_NET244_XI39/MM3059_g N_VSS_XI39/MM3059_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2391 XI39/NET10658 N_NET375_XI39/MM2391_g N_VSS_XI39/MM2391_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2380 N_NET476_XI39/MM2380_d N_NET376_XI39/MM2380_g N_VSS_XI39/MM2380_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2412 XI39/NET11222 N_NET377_XI39/MM2412_g N_VSS_XI39/MM2412_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2419 N_NET476_XI39/MM2419_d N_NET378_XI39/MM2419_g N_VSS_XI39/MM2419_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2348 XI39/NET10830 N_NET379_XI39/MM2348_g N_VSS_XI39/MM2348_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2355 N_NET476_XI39/MM2355_d N_NET380_XI39/MM2355_g N_VSS_XI39/MM2355_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2333 XI39/NET10890 N_NET381_XI39/MM2333_g N_VSS_XI39/MM2333_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2316 N_NET476_XI39/MM2316_d N_NET382_XI39/MM2316_g N_VSS_XI39/MM2316_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2478 XI39/NET11534 N_NET383_XI39/MM2478_g N_VSS_XI39/MM2478_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2483 N_NET476_XI39/MM2483_d N_NET384_XI39/MM2483_g N_VSS_XI39/MM2483_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2461 XI39/NET11026 N_NET385_XI39/MM2461_g N_VSS_XI39/MM2461_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2444 N_NET476_XI39/MM2444_d N_NET256_XI39/MM2444_g N_VSS_XI39/MM2444_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2525 XI39/NET11346 N_NET387_XI39/MM2525_g N_VSS_XI39/MM2525_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2508 N_NET476_XI39/MM2508_d N_NET388_XI39/MM2508_g N_VSS_XI39/MM2508_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2534 XI39/NET11310 N_NET389_XI39/MM2534_g N_VSS_XI39/MM2534_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2547 N_NET476_XI39/MM2547_d N_NET390_XI39/MM2547_g N_VSS_XI39/MM2547_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2220 XI39/NET10470 N_NET391_XI39/MM2220_g N_VSS_XI39/MM2220_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2227 N_NET476_XI39/MM2227_d N_NET262_XI39/MM2227_g N_VSS_XI39/MM2227_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2205 XI39/NET10530 N_NET263_XI39/MM2205_g N_VSS_XI39/MM2205_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2188 N_NET476_XI39/MM2188_d N_NET264_XI39/MM2188_g N_VSS_XI39/MM2188_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2269 XI39/NET10282 N_NET265_XI39/MM2269_g N_VSS_XI39/MM2269_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2252 N_NET476_XI39/MM2252_d N_NET396_XI39/MM2252_g N_VSS_XI39/MM2252_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2284 XI39/NET10222 N_NET267_XI39/MM2284_g N_VSS_XI39/MM2284_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2291 N_NET476_XI39/MM2291_d N_NET268_XI39/MM2291_g N_VSS_XI39/MM2291_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2137 XI39/NET9782 N_NET269_XI39/MM2137_g N_VSS_XI39/MM2137_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2124 N_NET476_XI39/MM2124_d N_NET270_XI39/MM2124_g N_VSS_XI39/MM2124_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2156 XI39/NET9706 N_NET401_XI39/MM2156_g N_VSS_XI39/MM2156_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2163 N_NET476_XI39/MM2163_d N_NET272_XI39/MM2163_g N_VSS_XI39/MM2163_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2092 XI39/NET9958 N_NET273_XI39/MM2092_g N_VSS_XI39/MM2092_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2099 N_NET476_XI39/MM2099_d N_NET404_XI39/MM2099_g N_VSS_XI39/MM2099_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2067 XI39/NET10018 N_NET405_XI39/MM2067_g N_VSS_XI39/MM2067_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3 N_NET476_XI39/MM3_d N_NET0390_XI39/MM3_g N_VSS_XI39/MM3_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3411 N_NET414_XI39/MM3411_d N_NET0133_XI39/MM3411_g N_VSS_XI39/MM3411_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3395 XI39/NET5642 N_NET280_XI39/MM3395_g N_VSS_XI39/MM3395_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3434 N_NET414_XI39/MM3434_d N_NET281_XI39/MM3434_g N_VSS_XI39/MM3434_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3441 XI39/NET5458 N_NET282_XI39/MM3441_g N_VSS_XI39/MM3441_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3371 N_NET414_XI39/MM3371_d N_NET153_XI39/MM3371_g N_VSS_XI39/MM3371_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3378 XI39/NET5710 N_NET284_XI39/MM3378_g N_VSS_XI39/MM3378_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3348 N_NET414_XI39/MM3348_d N_NET285_XI39/MM3348_g N_VSS_XI39/MM3348_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3341 XI39/NET3558 N_NET286_XI39/MM3341_g N_VSS_XI39/MM3341_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3498 N_NET414_XI39/MM3498_d N_NET287_XI39/MM3498_g N_VSS_XI39/MM3498_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3505 XI39/NET5202 N_NET158_XI39/MM3505_g N_VSS_XI39/MM3505_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3475 N_NET414_XI39/MM3475_d N_NET159_XI39/MM3475_g N_VSS_XI39/MM3475_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3458 XI39/NET5390 N_NET160_XI39/MM3458_g N_VSS_XI39/MM3458_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3539 N_NET414_XI39/MM3539_d N_NET291_XI39/MM3539_g N_VSS_XI39/MM3539_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3522 XI39/NET5134 N_NET162_XI39/MM3522_g N_VSS_XI39/MM3522_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3562 N_NET414_XI39/MM3562_d N_NET293_XI39/MM3562_g N_VSS_XI39/MM3562_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3569 XI39/NET4946 N_NET294_XI39/MM3569_g N_VSS_XI39/MM3569_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3243 N_NET414_XI39/MM3243_d N_NET295_XI39/MM3243_g N_VSS_XI39/MM3243_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3250 XI39/NET3922 N_NET296_XI39/MM3250_g N_VSS_XI39/MM3250_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3220 N_NET414_XI39/MM3220_d N_NET297_XI39/MM3220_g N_VSS_XI39/MM3220_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3203 XI39/NET4110 N_NET298_XI39/MM3203_g N_VSS_XI39/MM3203_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3284 N_NET414_XI39/MM3284_d N_NET299_XI39/MM3284_g N_VSS_XI39/MM3284_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3267 XI39/NET3854 N_NET170_XI39/MM3267_g N_VSS_XI39/MM3267_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3307 N_NET414_XI39/MM3307_d N_NET171_XI39/MM3307_g N_VSS_XI39/MM3307_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3314 XI39/NET3666 N_NET172_XI39/MM3314_g N_VSS_XI39/MM3314_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3156 N_NET414_XI39/MM3156_d N_NET303_XI39/MM3156_g N_VSS_XI39/MM3156_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3139 XI39/NET4366 N_NET304_XI39/MM3139_g N_VSS_XI39/MM3139_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3179 N_NET414_XI39/MM3179_d N_NET305_XI39/MM3179_g N_VSS_XI39/MM3179_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3186 XI39/NET4178 N_NET306_XI39/MM3186_g N_VSS_XI39/MM3186_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3115 N_NET414_XI39/MM3115_d N_NET307_XI39/MM3115_g N_VSS_XI39/MM3115_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3122 XI39/NET4434 N_NET308_XI39/MM3122_g N_VSS_XI39/MM3122_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3092 N_NET414_XI39/MM3092_d N_NET309_XI39/MM3092_g N_VSS_XI39/MM3092_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3075 XI39/NET4622 N_NET310_XI39/MM3075_g N_VSS_XI39/MM3075_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3844 N_NET414_XI39/MM3844_d N_NET311_XI39/MM3844_g N_VSS_XI39/MM3844_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3851 XI39/NET6118 N_NET312_XI39/MM3851_g N_VSS_XI39/MM3851_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3983 N_NET414_XI39/MM3983_d N_NET313_XI39/MM3983_g N_VSS_XI39/MM3983_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3966 XI39/NET7454 N_NET314_XI39/MM3966_g N_VSS_XI39/MM3966_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3885 N_NET414_XI39/MM3885_d N_NET315_XI39/MM3885_g N_VSS_XI39/MM3885_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3868 XI39/NET6050 N_NET316_XI39/MM3868_g N_VSS_XI39/MM3868_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3908 N_NET414_XI39/MM3908_d N_NET317_XI39/MM3908_g N_VSS_XI39/MM3908_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3915 XI39/NET5862 N_NET318_XI39/MM3915_g N_VSS_XI39/MM3915_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4063 N_NET414_XI39/MM4063_d N_NET319_XI39/MM4063_g N_VSS_XI39/MM4063_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4046 XI39/NET7134 N_NET320_XI39/MM4046_g N_VSS_XI39/MM4046_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3942 N_NET414_XI39/MM3942_d N_NET321_XI39/MM3942_g N_VSS_XI39/MM3942_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3949 XI39/NET7522 N_NET192_XI39/MM3949_g N_VSS_XI39/MM3949_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4022 N_NET414_XI39/MM4022_d N_NET193_XI39/MM4022_g N_VSS_XI39/MM4022_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4029 XI39/NET7202 N_NET194_XI39/MM4029_g N_VSS_XI39/MM4029_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4093 N_NET414_XI39/MM4093_d N_NET195_XI39/MM4093_g N_VSS_XI39/MM4093_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4076 XI39/NET7014 N_NET196_XI39/MM4076_g N_VSS_XI39/MM4076_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3795 N_NET414_XI39/MM3795_d N_NET197_XI39/MM3795_g N_VSS_XI39/MM3795_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3778 XI39/NET6410 N_NET198_XI39/MM3778_g N_VSS_XI39/MM3778_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3818 N_NET414_XI39/MM3818_d N_NET199_XI39/MM3818_g N_VSS_XI39/MM3818_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3825 XI39/NET6222 N_NET200_XI39/MM3825_g N_VSS_XI39/MM3825_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3754 N_NET414_XI39/MM3754_d N_NET331_XI39/MM3754_g N_VSS_XI39/MM3754_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3761 XI39/NET6478 N_NET332_XI39/MM3761_g N_VSS_XI39/MM3761_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3731 N_NET414_XI39/MM3731_d N_NET203_XI39/MM3731_g N_VSS_XI39/MM3731_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3714 XI39/NET6666 N_NET204_XI39/MM3714_g N_VSS_XI39/MM3714_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3626 N_NET414_XI39/MM3626_d N_NET205_XI39/MM3626_g N_VSS_XI39/MM3626_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3633 XI39/NET4690 N_NET206_XI39/MM3633_g N_VSS_XI39/MM3633_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3603 N_NET414_XI39/MM3603_d N_NET207_XI39/MM3603_g N_VSS_XI39/MM3603_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3586 XI39/NET4878 N_NET338_XI39/MM3586_g N_VSS_XI39/MM3586_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3667 N_NET414_XI39/MM3667_d N_NET339_XI39/MM3667_g N_VSS_XI39/MM3667_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3650 XI39/NET6922 N_NET340_XI39/MM3650_g N_VSS_XI39/MM3650_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3683 N_NET414_XI39/MM3683_d N_NET211_XI39/MM3683_g N_VSS_XI39/MM3683_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3690 XI39/NET6762 N_NET212_XI39/MM3690_g N_VSS_XI39/MM3690_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2731 N_NET414_XI39/MM2731_d N_NET214_XI39/MM2731_g N_VSS_XI39/MM2731_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2738 XI39/NET8914 N_NET215_XI39/MM2738_g N_VSS_XI39/MM2738_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2708 N_NET414_XI39/MM2708_d N_NET216_XI39/MM2708_g N_VSS_XI39/MM2708_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2691 XI39/NET9098 N_NET346_XI39/MM2691_g N_VSS_XI39/MM2691_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2772 N_NET414_XI39/MM2772_d N_NET347_XI39/MM2772_g N_VSS_XI39/MM2772_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2755 XI39/NET8846 N_NET348_XI39/MM2755_g N_VSS_XI39/MM2755_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2795 N_NET414_XI39/MM2795_d N_NET349_XI39/MM2795_g N_VSS_XI39/MM2795_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2802 XI39/NET8658 N_NET350_XI39/MM2802_g N_VSS_XI39/MM2802_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2644 N_NET414_XI39/MM2644_d N_NET351_XI39/MM2644_g N_VSS_XI39/MM2644_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2627 XI39/NET9354 N_NET352_XI39/MM2627_g N_VSS_XI39/MM2627_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2667 N_NET414_XI39/MM2667_d N_NET224_XI39/MM2667_g N_VSS_XI39/MM2667_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2674 XI39/NET9166 N_NET225_XI39/MM2674_g N_VSS_XI39/MM2674_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2603 N_NET414_XI39/MM2603_d N_NET226_XI39/MM2603_g N_VSS_XI39/MM2603_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2610 XI39/NET9422 N_NET356_XI39/MM2610_g N_VSS_XI39/MM2610_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2580 N_NET414_XI39/MM2580_d N_NET357_XI39/MM2580_g N_VSS_XI39/MM2580_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2563 XI39/NET9610 N_NET358_XI39/MM2563_g N_VSS_XI39/MM2563_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2900 N_NET414_XI39/MM2900_d N_NET230_XI39/MM2900_g N_VSS_XI39/MM2900_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2883 XI39/NET8334 N_NET360_XI39/MM2883_g N_VSS_XI39/MM2883_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2923 N_NET414_XI39/MM2923_d N_NET361_XI39/MM2923_g N_VSS_XI39/MM2923_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2930 XI39/NET8146 N_NET233_XI39/MM2930_g N_VSS_XI39/MM2930_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2859 N_NET414_XI39/MM2859_d N_NET234_XI39/MM2859_g N_VSS_XI39/MM2859_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2866 XI39/NET8402 N_NET235_XI39/MM2866_g N_VSS_XI39/MM2866_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2836 N_NET414_XI39/MM2836_d N_NET365_XI39/MM2836_g N_VSS_XI39/MM2836_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2819 XI39/NET8590 N_NET366_XI39/MM2819_g N_VSS_XI39/MM2819_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2987 N_NET414_XI39/MM2987_d N_NET367_XI39/MM2987_g N_VSS_XI39/MM2987_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2994 XI39/NET7890 N_NET368_XI39/MM2994_g N_VSS_XI39/MM2994_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2964 N_NET414_XI39/MM2964_d N_NET369_XI39/MM2964_g N_VSS_XI39/MM2964_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2947 XI39/NET8078 N_NET370_XI39/MM2947_g N_VSS_XI39/MM2947_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3028 N_NET414_XI39/MM3028_d N_NET371_XI39/MM3028_g N_VSS_XI39/MM3028_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3011 XI39/NET7822 N_NET242_XI39/MM3011_g N_VSS_XI39/MM3011_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3051 N_NET414_XI39/MM3051_d N_NET373_XI39/MM3051_g N_VSS_XI39/MM3051_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3058 XI39/NET7634 N_NET244_XI39/MM3058_g N_VSS_XI39/MM3058_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2388 N_NET414_XI39/MM2388_d N_NET375_XI39/MM2388_g N_VSS_XI39/MM2388_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2371 XI39/NET10738 N_NET376_XI39/MM2371_g N_VSS_XI39/MM2371_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2411 N_NET414_XI39/MM2411_d N_NET377_XI39/MM2411_g N_VSS_XI39/MM2411_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2418 XI39/NET11198 N_NET378_XI39/MM2418_g N_VSS_XI39/MM2418_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2347 N_NET414_XI39/MM2347_d N_NET379_XI39/MM2347_g N_VSS_XI39/MM2347_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2354 XI39/NET10806 N_NET380_XI39/MM2354_g N_VSS_XI39/MM2354_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2324 N_NET414_XI39/MM2324_d N_NET381_XI39/MM2324_g N_VSS_XI39/MM2324_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2307 XI39/NET10994 N_NET382_XI39/MM2307_g N_VSS_XI39/MM2307_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2475 N_NET414_XI39/MM2475_d N_NET383_XI39/MM2475_g N_VSS_XI39/MM2475_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2482 XI39/NET11518 N_NET384_XI39/MM2482_g N_VSS_XI39/MM2482_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2452 N_NET414_XI39/MM2452_d N_NET385_XI39/MM2452_g N_VSS_XI39/MM2452_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2435 XI39/NET11130 N_NET256_XI39/MM2435_g N_VSS_XI39/MM2435_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2516 N_NET414_XI39/MM2516_d N_NET387_XI39/MM2516_g N_VSS_XI39/MM2516_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2499 XI39/NET11450 N_NET388_XI39/MM2499_g N_VSS_XI39/MM2499_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2539 N_NET414_XI39/MM2539_d N_NET389_XI39/MM2539_g N_VSS_XI39/MM2539_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2546 XI39/NET11638 N_NET390_XI39/MM2546_g N_VSS_XI39/MM2546_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2219 N_NET414_XI39/MM2219_d N_NET391_XI39/MM2219_g N_VSS_XI39/MM2219_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2226 XI39/NET10450 N_NET262_XI39/MM2226_g N_VSS_XI39/MM2226_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2196 N_NET414_XI39/MM2196_d N_NET263_XI39/MM2196_g N_VSS_XI39/MM2196_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2179 XI39/NET10630 N_NET264_XI39/MM2179_g N_VSS_XI39/MM2179_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2260 N_NET414_XI39/MM2260_d N_NET265_XI39/MM2260_g N_VSS_XI39/MM2260_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2243 XI39/NET10382 N_NET396_XI39/MM2243_g N_VSS_XI39/MM2243_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2283 N_NET414_XI39/MM2283_d N_NET267_XI39/MM2283_g N_VSS_XI39/MM2283_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2290 XI39/NET10202 N_NET268_XI39/MM2290_g N_VSS_XI39/MM2290_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2132 N_NET414_XI39/MM2132_d N_NET269_XI39/MM2132_g N_VSS_XI39/MM2132_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2115 XI39/NET9866 N_NET270_XI39/MM2115_g N_VSS_XI39/MM2115_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2155 N_NET414_XI39/MM2155_d N_NET401_XI39/MM2155_g N_VSS_XI39/MM2155_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2162 XI39/NET9686 N_NET272_XI39/MM2162_g N_VSS_XI39/MM2162_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2091 N_NET414_XI39/MM2091_d N_NET273_XI39/MM2091_g N_VSS_XI39/MM2091_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2098 XI39/NET9938 N_NET404_XI39/MM2098_g N_VSS_XI39/MM2098_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2068 N_NET414_XI39/MM2068_d N_NET405_XI39/MM2068_g N_VSS_XI39/MM2068_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM12 XI39/NET10090 N_NET0390_XI39/MM12_g N_VSS_XI39/MM12_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI29/XI0/MM43 N_NET414_XI29/XI0/MM43_d N_XI29/XI0/NET211_XI29/XI0/MM43_g
+ N_NET064_XI29/XI0/MM43_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI29/XI0/XI12/MM1 N_XI29/XI0/NET211_XI29/XI0/XI12/MM1_d
+ N_NET466_XI29/XI0/XI12/MM1_g N_VSS_XI29/XI0/XI12/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI29/XI0/MM44 N_NET415_XI29/XI0/MM44_d N_XI29/XI0/NET203_XI29/XI0/MM44_g
+ N_NET064_XI29/XI0/MM44_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI29/XI0/XI13/MM1 N_XI29/XI0/NET203_XI29/XI0/XI13/MM1_d
+ N_NET465_XI29/XI0/XI13/MM1_g N_VSS_XI29/XI0/XI13/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI39/MM3410 XI39/NET5582 N_NET0133_XI39/MM3410_g N_VSS_XI39/MM3410_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3402 N_NET415_XI39/MM3402_d N_NET280_XI39/MM3402_g N_VSS_XI39/MM3402_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3425 XI39/NET5522 N_NET281_XI39/MM3425_g N_VSS_XI39/MM3425_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3444 N_NET415_XI39/MM3444_d N_NET282_XI39/MM3444_g N_VSS_XI39/MM3444_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3362 XI39/NET5774 N_NET153_XI39/MM3362_g N_VSS_XI39/MM3362_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3381 N_NET415_XI39/MM3381_d N_NET284_XI39/MM3381_g N_VSS_XI39/MM3381_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3347 XI39/NET3534 N_NET285_XI39/MM3347_g N_VSS_XI39/MM3347_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3338 N_NET415_XI39/MM3338_d N_NET286_XI39/MM3338_g N_VSS_XI39/MM3338_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3489 XI39/NET5266 N_NET287_XI39/MM3489_g N_VSS_XI39/MM3489_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3508 N_NET415_XI39/MM3508_d N_NET158_XI39/MM3508_g N_VSS_XI39/MM3508_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3474 XI39/NET5326 N_NET159_XI39/MM3474_g N_VSS_XI39/MM3474_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3465 N_NET415_XI39/MM3465_d N_NET160_XI39/MM3465_g N_VSS_XI39/MM3465_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3538 XI39/NET5070 N_NET291_XI39/MM3538_g N_VSS_XI39/MM3538_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3529 N_NET415_XI39/MM3529_d N_NET162_XI39/MM3529_g N_VSS_XI39/MM3529_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3553 XI39/NET5010 N_NET293_XI39/MM3553_g N_VSS_XI39/MM3553_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3572 N_NET415_XI39/MM3572_d N_NET294_XI39/MM3572_g N_VSS_XI39/MM3572_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3234 XI39/NET3986 N_NET295_XI39/MM3234_g N_VSS_XI39/MM3234_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3253 N_NET415_XI39/MM3253_d N_NET296_XI39/MM3253_g N_VSS_XI39/MM3253_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3219 XI39/NET4046 N_NET297_XI39/MM3219_g N_VSS_XI39/MM3219_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3210 N_NET415_XI39/MM3210_d N_NET298_XI39/MM3210_g N_VSS_XI39/MM3210_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3283 XI39/NET3790 N_NET299_XI39/MM3283_g N_VSS_XI39/MM3283_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3274 N_NET415_XI39/MM3274_d N_NET170_XI39/MM3274_g N_VSS_XI39/MM3274_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3298 XI39/NET3730 N_NET171_XI39/MM3298_g N_VSS_XI39/MM3298_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3317 N_NET415_XI39/MM3317_d N_NET172_XI39/MM3317_g N_VSS_XI39/MM3317_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3155 XI39/NET4302 N_NET303_XI39/MM3155_g N_VSS_XI39/MM3155_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3146 N_NET415_XI39/MM3146_d N_NET304_XI39/MM3146_g N_VSS_XI39/MM3146_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3170 XI39/NET4242 N_NET305_XI39/MM3170_g N_VSS_XI39/MM3170_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3189 N_NET415_XI39/MM3189_d N_NET306_XI39/MM3189_g N_VSS_XI39/MM3189_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3106 XI39/NET4498 N_NET307_XI39/MM3106_g N_VSS_XI39/MM3106_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3125 N_NET415_XI39/MM3125_d N_NET308_XI39/MM3125_g N_VSS_XI39/MM3125_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3091 XI39/NET4558 N_NET309_XI39/MM3091_g N_VSS_XI39/MM3091_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3082 N_NET415_XI39/MM3082_d N_NET310_XI39/MM3082_g N_VSS_XI39/MM3082_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3997 XI39/NET7330 N_NET311_XI39/MM3997_g N_VSS_XI39/MM3997_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3854 N_NET415_XI39/MM3854_d N_NET312_XI39/MM3854_g N_VSS_XI39/MM3854_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3982 XI39/NET7390 N_NET313_XI39/MM3982_g N_VSS_XI39/MM3982_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3973 N_NET415_XI39/MM3973_d N_NET314_XI39/MM3973_g N_VSS_XI39/MM3973_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3884 XI39/NET5986 N_NET315_XI39/MM3884_g N_VSS_XI39/MM3884_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3875 N_NET415_XI39/MM3875_d N_NET316_XI39/MM3875_g N_VSS_XI39/MM3875_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3899 XI39/NET5926 N_NET317_XI39/MM3899_g N_VSS_XI39/MM3899_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3918 N_NET415_XI39/MM3918_d N_NET318_XI39/MM3918_g N_VSS_XI39/MM3918_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4062 XI39/NET7070 N_NET319_XI39/MM4062_g N_VSS_XI39/MM4062_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4053 N_NET415_XI39/MM4053_d N_NET320_XI39/MM4053_g N_VSS_XI39/MM4053_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3937 XI39/NET7570 N_NET321_XI39/MM3937_g N_VSS_XI39/MM3937_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3952 N_NET415_XI39/MM3952_d N_NET192_XI39/MM3952_g N_VSS_XI39/MM3952_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4013 XI39/NET7266 N_NET193_XI39/MM4013_g N_VSS_XI39/MM4013_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4032 N_NET415_XI39/MM4032_d N_NET194_XI39/MM4032_g N_VSS_XI39/MM4032_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4004 XI39/NET7302 N_NET195_XI39/MM4004_g N_VSS_XI39/MM4004_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4083 N_NET415_XI39/MM4083_d N_NET196_XI39/MM4083_g N_VSS_XI39/MM4083_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3794 XI39/NET6346 N_NET197_XI39/MM3794_g N_VSS_XI39/MM3794_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3785 N_NET415_XI39/MM3785_d N_NET198_XI39/MM3785_g N_VSS_XI39/MM3785_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3809 XI39/NET6286 N_NET199_XI39/MM3809_g N_VSS_XI39/MM3809_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3828 N_NET415_XI39/MM3828_d N_NET200_XI39/MM3828_g N_VSS_XI39/MM3828_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3745 XI39/NET6542 N_NET331_XI39/MM3745_g N_VSS_XI39/MM3745_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3764 N_NET415_XI39/MM3764_d N_NET332_XI39/MM3764_g N_VSS_XI39/MM3764_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3730 XI39/NET6602 N_NET203_XI39/MM3730_g N_VSS_XI39/MM3730_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3721 N_NET415_XI39/MM3721_d N_NET204_XI39/MM3721_g N_VSS_XI39/MM3721_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3617 XI39/NET4754 N_NET205_XI39/MM3617_g N_VSS_XI39/MM3617_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3636 N_NET415_XI39/MM3636_d N_NET206_XI39/MM3636_g N_VSS_XI39/MM3636_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3602 XI39/NET4814 N_NET207_XI39/MM3602_g N_VSS_XI39/MM3602_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3593 N_NET415_XI39/MM3593_d N_NET338_XI39/MM3593_g N_VSS_XI39/MM3593_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3666 XI39/NET6858 N_NET339_XI39/MM3666_g N_VSS_XI39/MM3666_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3657 N_NET415_XI39/MM3657_d N_NET340_XI39/MM3657_g N_VSS_XI39/MM3657_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3682 XI39/NET6794 N_NET211_XI39/MM3682_g N_VSS_XI39/MM3682_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3693 N_NET415_XI39/MM3693_d N_NET212_XI39/MM3693_g N_VSS_XI39/MM3693_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2722 XI39/NET8974 N_NET214_XI39/MM2722_g N_VSS_XI39/MM2722_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2741 N_NET415_XI39/MM2741_d N_NET215_XI39/MM2741_g N_VSS_XI39/MM2741_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2707 XI39/NET9034 N_NET216_XI39/MM2707_g N_VSS_XI39/MM2707_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2698 N_NET415_XI39/MM2698_d N_NET346_XI39/MM2698_g N_VSS_XI39/MM2698_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2771 XI39/NET8782 N_NET347_XI39/MM2771_g N_VSS_XI39/MM2771_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2762 N_NET415_XI39/MM2762_d N_NET348_XI39/MM2762_g N_VSS_XI39/MM2762_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2786 XI39/NET8722 N_NET349_XI39/MM2786_g N_VSS_XI39/MM2786_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2805 N_NET415_XI39/MM2805_d N_NET350_XI39/MM2805_g N_VSS_XI39/MM2805_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2643 XI39/NET9290 N_NET351_XI39/MM2643_g N_VSS_XI39/MM2643_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2634 N_NET415_XI39/MM2634_d N_NET352_XI39/MM2634_g N_VSS_XI39/MM2634_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2658 XI39/NET9230 N_NET224_XI39/MM2658_g N_VSS_XI39/MM2658_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2677 N_NET415_XI39/MM2677_d N_NET225_XI39/MM2677_g N_VSS_XI39/MM2677_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2594 XI39/NET9486 N_NET226_XI39/MM2594_g N_VSS_XI39/MM2594_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2613 N_NET415_XI39/MM2613_d N_NET356_XI39/MM2613_g N_VSS_XI39/MM2613_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2579 XI39/NET9546 N_NET357_XI39/MM2579_g N_VSS_XI39/MM2579_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2570 N_NET415_XI39/MM2570_d N_NET358_XI39/MM2570_g N_VSS_XI39/MM2570_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2899 XI39/NET8270 N_NET230_XI39/MM2899_g N_VSS_XI39/MM2899_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2890 N_NET415_XI39/MM2890_d N_NET360_XI39/MM2890_g N_VSS_XI39/MM2890_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2914 XI39/NET8210 N_NET361_XI39/MM2914_g N_VSS_XI39/MM2914_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2933 N_NET415_XI39/MM2933_d N_NET233_XI39/MM2933_g N_VSS_XI39/MM2933_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2850 XI39/NET8466 N_NET234_XI39/MM2850_g N_VSS_XI39/MM2850_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2869 N_NET415_XI39/MM2869_d N_NET235_XI39/MM2869_g N_VSS_XI39/MM2869_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2835 XI39/NET8526 N_NET365_XI39/MM2835_g N_VSS_XI39/MM2835_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2826 N_NET415_XI39/MM2826_d N_NET366_XI39/MM2826_g N_VSS_XI39/MM2826_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2978 XI39/NET7954 N_NET367_XI39/MM2978_g N_VSS_XI39/MM2978_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2997 N_NET415_XI39/MM2997_d N_NET368_XI39/MM2997_g N_VSS_XI39/MM2997_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2963 XI39/NET8014 N_NET369_XI39/MM2963_g N_VSS_XI39/MM2963_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2954 N_NET415_XI39/MM2954_d N_NET370_XI39/MM2954_g N_VSS_XI39/MM2954_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3027 XI39/NET7758 N_NET371_XI39/MM3027_g N_VSS_XI39/MM3027_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3018 N_NET415_XI39/MM3018_d N_NET242_XI39/MM3018_g N_VSS_XI39/MM3018_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3042 XI39/NET7698 N_NET373_XI39/MM3042_g N_VSS_XI39/MM3042_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3061 N_NET415_XI39/MM3061_d N_NET244_XI39/MM3061_g N_VSS_XI39/MM3061_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2397 XI39/NET11282 N_NET375_XI39/MM2397_g N_VSS_XI39/MM2397_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2378 N_NET415_XI39/MM2378_d N_NET376_XI39/MM2378_g N_VSS_XI39/MM2378_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2402 XI39/NET11262 N_NET377_XI39/MM2402_g N_VSS_XI39/MM2402_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2421 N_NET415_XI39/MM2421_d N_NET378_XI39/MM2421_g N_VSS_XI39/MM2421_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2338 XI39/NET10870 N_NET379_XI39/MM2338_g N_VSS_XI39/MM2338_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2357 N_NET415_XI39/MM2357_d N_NET380_XI39/MM2357_g N_VSS_XI39/MM2357_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2323 XI39/NET10930 N_NET381_XI39/MM2323_g N_VSS_XI39/MM2323_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2314 N_NET415_XI39/MM2314_d N_NET382_XI39/MM2314_g N_VSS_XI39/MM2314_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2468 XI39/NET11574 N_NET383_XI39/MM2468_g N_VSS_XI39/MM2468_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2485 N_NET415_XI39/MM2485_d N_NET384_XI39/MM2485_g N_VSS_XI39/MM2485_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2451 XI39/NET11066 N_NET385_XI39/MM2451_g N_VSS_XI39/MM2451_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2442 N_NET415_XI39/MM2442_d N_NET256_XI39/MM2442_g N_VSS_XI39/MM2442_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2515 XI39/NET11386 N_NET387_XI39/MM2515_g N_VSS_XI39/MM2515_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2506 N_NET415_XI39/MM2506_d N_NET388_XI39/MM2506_g N_VSS_XI39/MM2506_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2540 XI39/NET11662 N_NET389_XI39/MM2540_g N_VSS_XI39/MM2540_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2549 N_NET415_XI39/MM2549_d N_NET390_XI39/MM2549_g N_VSS_XI39/MM2549_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2210 XI39/NET10510 N_NET391_XI39/MM2210_g N_VSS_XI39/MM2210_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2229 N_NET415_XI39/MM2229_d N_NET262_XI39/MM2229_g N_VSS_XI39/MM2229_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2195 XI39/NET10570 N_NET263_XI39/MM2195_g N_VSS_XI39/MM2195_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2186 N_NET415_XI39/MM2186_d N_NET264_XI39/MM2186_g N_VSS_XI39/MM2186_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2259 XI39/NET10322 N_NET265_XI39/MM2259_g N_VSS_XI39/MM2259_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2250 N_NET415_XI39/MM2250_d N_NET396_XI39/MM2250_g N_VSS_XI39/MM2250_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2274 XI39/NET10262 N_NET267_XI39/MM2274_g N_VSS_XI39/MM2274_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2293 N_NET415_XI39/MM2293_d N_NET268_XI39/MM2293_g N_VSS_XI39/MM2293_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2131 XI39/NET9806 N_NET269_XI39/MM2131_g N_VSS_XI39/MM2131_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2122 N_NET415_XI39/MM2122_d N_NET270_XI39/MM2122_g N_VSS_XI39/MM2122_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2146 XI39/NET9746 N_NET401_XI39/MM2146_g N_VSS_XI39/MM2146_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2165 N_NET415_XI39/MM2165_d N_NET272_XI39/MM2165_g N_VSS_XI39/MM2165_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2082 XI39/NET9998 N_NET273_XI39/MM2082_g N_VSS_XI39/MM2082_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2101 N_NET415_XI39/MM2101_d N_NET404_XI39/MM2101_g N_VSS_XI39/MM2101_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2077 XI39/NET10122 N_NET405_XI39/MM2077_g N_VSS_XI39/MM2077_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM5 N_NET415_XI39/MM5_d N_NET0390_XI39/MM5_g N_VSS_XI39/MM5_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI29/XI0/MM45 N_NET416_XI29/XI0/MM45_d N_XI29/XI0/NET219_XI29/XI0/MM45_g
+ N_NET064_XI29/XI0/MM45_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI29/XI0/XI14/MM1 N_XI29/XI0/NET219_XI29/XI0/XI14/MM1_d
+ N_NET464_XI29/XI0/XI14/MM1_g N_VSS_XI29/XI0/XI14/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI29/XI0/MM46 N_NET417_XI29/XI0/MM46_d N_XI29/XI0/NET207_XI29/XI0/MM46_g
+ N_NET064_XI29/XI0/MM46_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI29/XI0/XI15/MM1 N_XI29/XI0/NET207_XI29/XI0/XI15/MM1_d
+ N_NET463_XI29/XI0/XI15/MM1_g N_VSS_XI29/XI0/XI15/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI39/MM3413 N_NET416_XI39/MM3413_d N_NET0133_XI39/MM3413_g N_VSS_XI39/MM3413_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3397 XI39/NET5634 N_NET280_XI39/MM3397_g N_VSS_XI39/MM3397_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3432 N_NET416_XI39/MM3432_d N_NET281_XI39/MM3432_g N_VSS_XI39/MM3432_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3443 XI39/NET5450 N_NET282_XI39/MM3443_g N_VSS_XI39/MM3443_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3369 N_NET416_XI39/MM3369_d N_NET153_XI39/MM3369_g N_VSS_XI39/MM3369_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3380 XI39/NET5702 N_NET284_XI39/MM3380_g N_VSS_XI39/MM3380_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3350 N_NET416_XI39/MM3350_d N_NET285_XI39/MM3350_g N_VSS_XI39/MM3350_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3335 XI39/NET3582 N_NET286_XI39/MM3335_g N_VSS_XI39/MM3335_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3496 N_NET416_XI39/MM3496_d N_NET287_XI39/MM3496_g N_VSS_XI39/MM3496_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3507 XI39/NET5194 N_NET158_XI39/MM3507_g N_VSS_XI39/MM3507_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3477 N_NET416_XI39/MM3477_d N_NET159_XI39/MM3477_g N_VSS_XI39/MM3477_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3460 XI39/NET5382 N_NET160_XI39/MM3460_g N_VSS_XI39/MM3460_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3541 N_NET416_XI39/MM3541_d N_NET291_XI39/MM3541_g N_VSS_XI39/MM3541_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3524 XI39/NET5126 N_NET162_XI39/MM3524_g N_VSS_XI39/MM3524_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3560 N_NET416_XI39/MM3560_d N_NET293_XI39/MM3560_g N_VSS_XI39/MM3560_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3571 XI39/NET4938 N_NET294_XI39/MM3571_g N_VSS_XI39/MM3571_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3241 N_NET416_XI39/MM3241_d N_NET295_XI39/MM3241_g N_VSS_XI39/MM3241_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3252 XI39/NET3914 N_NET296_XI39/MM3252_g N_VSS_XI39/MM3252_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3222 N_NET416_XI39/MM3222_d N_NET297_XI39/MM3222_g N_VSS_XI39/MM3222_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3205 XI39/NET4102 N_NET298_XI39/MM3205_g N_VSS_XI39/MM3205_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3286 N_NET416_XI39/MM3286_d N_NET299_XI39/MM3286_g N_VSS_XI39/MM3286_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3269 XI39/NET3846 N_NET170_XI39/MM3269_g N_VSS_XI39/MM3269_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3305 N_NET416_XI39/MM3305_d N_NET171_XI39/MM3305_g N_VSS_XI39/MM3305_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3316 XI39/NET3658 N_NET172_XI39/MM3316_g N_VSS_XI39/MM3316_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3158 N_NET416_XI39/MM3158_d N_NET303_XI39/MM3158_g N_VSS_XI39/MM3158_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3141 XI39/NET4358 N_NET304_XI39/MM3141_g N_VSS_XI39/MM3141_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3177 N_NET416_XI39/MM3177_d N_NET305_XI39/MM3177_g N_VSS_XI39/MM3177_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3188 XI39/NET4170 N_NET306_XI39/MM3188_g N_VSS_XI39/MM3188_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3113 N_NET416_XI39/MM3113_d N_NET307_XI39/MM3113_g N_VSS_XI39/MM3113_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3124 XI39/NET4426 N_NET308_XI39/MM3124_g N_VSS_XI39/MM3124_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3094 N_NET416_XI39/MM3094_d N_NET309_XI39/MM3094_g N_VSS_XI39/MM3094_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3077 XI39/NET4614 N_NET310_XI39/MM3077_g N_VSS_XI39/MM3077_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3842 N_NET416_XI39/MM3842_d N_NET311_XI39/MM3842_g N_VSS_XI39/MM3842_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3853 XI39/NET6110 N_NET312_XI39/MM3853_g N_VSS_XI39/MM3853_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3985 N_NET416_XI39/MM3985_d N_NET313_XI39/MM3985_g N_VSS_XI39/MM3985_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3968 XI39/NET7446 N_NET314_XI39/MM3968_g N_VSS_XI39/MM3968_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3887 N_NET416_XI39/MM3887_d N_NET315_XI39/MM3887_g N_VSS_XI39/MM3887_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3870 XI39/NET6042 N_NET316_XI39/MM3870_g N_VSS_XI39/MM3870_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3906 N_NET416_XI39/MM3906_d N_NET317_XI39/MM3906_g N_VSS_XI39/MM3906_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3917 XI39/NET5854 N_NET318_XI39/MM3917_g N_VSS_XI39/MM3917_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4065 N_NET416_XI39/MM4065_d N_NET319_XI39/MM4065_g N_VSS_XI39/MM4065_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4048 XI39/NET7126 N_NET320_XI39/MM4048_g N_VSS_XI39/MM4048_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3940 N_NET416_XI39/MM3940_d N_NET321_XI39/MM3940_g N_VSS_XI39/MM3940_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3951 XI39/NET7514 N_NET192_XI39/MM3951_g N_VSS_XI39/MM3951_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4020 N_NET416_XI39/MM4020_d N_NET193_XI39/MM4020_g N_VSS_XI39/MM4020_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4031 XI39/NET7194 N_NET194_XI39/MM4031_g N_VSS_XI39/MM4031_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4001 N_NET416_XI39/MM4001_d N_NET195_XI39/MM4001_g N_VSS_XI39/MM4001_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4078 XI39/NET7006 N_NET196_XI39/MM4078_g N_VSS_XI39/MM4078_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3797 N_NET416_XI39/MM3797_d N_NET197_XI39/MM3797_g N_VSS_XI39/MM3797_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3780 XI39/NET6402 N_NET198_XI39/MM3780_g N_VSS_XI39/MM3780_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3816 N_NET416_XI39/MM3816_d N_NET199_XI39/MM3816_g N_VSS_XI39/MM3816_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3827 XI39/NET6214 N_NET200_XI39/MM3827_g N_VSS_XI39/MM3827_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3752 N_NET416_XI39/MM3752_d N_NET331_XI39/MM3752_g N_VSS_XI39/MM3752_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3763 XI39/NET6470 N_NET332_XI39/MM3763_g N_VSS_XI39/MM3763_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3733 N_NET416_XI39/MM3733_d N_NET203_XI39/MM3733_g N_VSS_XI39/MM3733_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3716 XI39/NET6658 N_NET204_XI39/MM3716_g N_VSS_XI39/MM3716_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3624 N_NET416_XI39/MM3624_d N_NET205_XI39/MM3624_g N_VSS_XI39/MM3624_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3635 XI39/NET4682 N_NET206_XI39/MM3635_g N_VSS_XI39/MM3635_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3605 N_NET416_XI39/MM3605_d N_NET207_XI39/MM3605_g N_VSS_XI39/MM3605_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3588 XI39/NET4870 N_NET338_XI39/MM3588_g N_VSS_XI39/MM3588_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3669 N_NET416_XI39/MM3669_d N_NET339_XI39/MM3669_g N_VSS_XI39/MM3669_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3652 XI39/NET6914 N_NET340_XI39/MM3652_g N_VSS_XI39/MM3652_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3685 N_NET416_XI39/MM3685_d N_NET211_XI39/MM3685_g N_VSS_XI39/MM3685_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3692 XI39/NET6754 N_NET212_XI39/MM3692_g N_VSS_XI39/MM3692_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2729 N_NET416_XI39/MM2729_d N_NET214_XI39/MM2729_g N_VSS_XI39/MM2729_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2740 XI39/NET8906 N_NET215_XI39/MM2740_g N_VSS_XI39/MM2740_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2710 N_NET416_XI39/MM2710_d N_NET216_XI39/MM2710_g N_VSS_XI39/MM2710_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2693 XI39/NET9090 N_NET346_XI39/MM2693_g N_VSS_XI39/MM2693_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2774 N_NET416_XI39/MM2774_d N_NET347_XI39/MM2774_g N_VSS_XI39/MM2774_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2757 XI39/NET8838 N_NET348_XI39/MM2757_g N_VSS_XI39/MM2757_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2793 N_NET416_XI39/MM2793_d N_NET349_XI39/MM2793_g N_VSS_XI39/MM2793_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2804 XI39/NET8650 N_NET350_XI39/MM2804_g N_VSS_XI39/MM2804_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2646 N_NET416_XI39/MM2646_d N_NET351_XI39/MM2646_g N_VSS_XI39/MM2646_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2629 XI39/NET9346 N_NET352_XI39/MM2629_g N_VSS_XI39/MM2629_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2665 N_NET416_XI39/MM2665_d N_NET224_XI39/MM2665_g N_VSS_XI39/MM2665_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2676 XI39/NET9158 N_NET225_XI39/MM2676_g N_VSS_XI39/MM2676_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2601 N_NET416_XI39/MM2601_d N_NET226_XI39/MM2601_g N_VSS_XI39/MM2601_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2612 XI39/NET9414 N_NET356_XI39/MM2612_g N_VSS_XI39/MM2612_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2582 N_NET416_XI39/MM2582_d N_NET357_XI39/MM2582_g N_VSS_XI39/MM2582_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2565 XI39/NET9602 N_NET358_XI39/MM2565_g N_VSS_XI39/MM2565_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2902 N_NET416_XI39/MM2902_d N_NET230_XI39/MM2902_g N_VSS_XI39/MM2902_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2885 XI39/NET8326 N_NET360_XI39/MM2885_g N_VSS_XI39/MM2885_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2921 N_NET416_XI39/MM2921_d N_NET361_XI39/MM2921_g N_VSS_XI39/MM2921_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2932 XI39/NET8138 N_NET233_XI39/MM2932_g N_VSS_XI39/MM2932_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2857 N_NET416_XI39/MM2857_d N_NET234_XI39/MM2857_g N_VSS_XI39/MM2857_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2868 XI39/NET8394 N_NET235_XI39/MM2868_g N_VSS_XI39/MM2868_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2838 N_NET416_XI39/MM2838_d N_NET365_XI39/MM2838_g N_VSS_XI39/MM2838_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2821 XI39/NET8582 N_NET366_XI39/MM2821_g N_VSS_XI39/MM2821_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2985 N_NET416_XI39/MM2985_d N_NET367_XI39/MM2985_g N_VSS_XI39/MM2985_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2996 XI39/NET7882 N_NET368_XI39/MM2996_g N_VSS_XI39/MM2996_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2966 N_NET416_XI39/MM2966_d N_NET369_XI39/MM2966_g N_VSS_XI39/MM2966_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2949 XI39/NET8070 N_NET370_XI39/MM2949_g N_VSS_XI39/MM2949_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3030 N_NET416_XI39/MM3030_d N_NET371_XI39/MM3030_g N_VSS_XI39/MM3030_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3013 XI39/NET7814 N_NET242_XI39/MM3013_g N_VSS_XI39/MM3013_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3049 N_NET416_XI39/MM3049_d N_NET373_XI39/MM3049_g N_VSS_XI39/MM3049_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3060 XI39/NET7626 N_NET244_XI39/MM3060_g N_VSS_XI39/MM3060_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2390 N_NET416_XI39/MM2390_d N_NET375_XI39/MM2390_g N_VSS_XI39/MM2390_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2373 XI39/NET10730 N_NET376_XI39/MM2373_g N_VSS_XI39/MM2373_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2409 N_NET416_XI39/MM2409_d N_NET377_XI39/MM2409_g N_VSS_XI39/MM2409_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2420 XI39/NET11190 N_NET378_XI39/MM2420_g N_VSS_XI39/MM2420_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2345 N_NET416_XI39/MM2345_d N_NET379_XI39/MM2345_g N_VSS_XI39/MM2345_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2356 XI39/NET10798 N_NET380_XI39/MM2356_g N_VSS_XI39/MM2356_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2326 N_NET416_XI39/MM2326_d N_NET381_XI39/MM2326_g N_VSS_XI39/MM2326_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2309 XI39/NET10986 N_NET382_XI39/MM2309_g N_VSS_XI39/MM2309_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2473 N_NET416_XI39/MM2473_d N_NET383_XI39/MM2473_g N_VSS_XI39/MM2473_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2484 XI39/NET11510 N_NET384_XI39/MM2484_g N_VSS_XI39/MM2484_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2454 N_NET416_XI39/MM2454_d N_NET385_XI39/MM2454_g N_VSS_XI39/MM2454_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2437 XI39/NET11122 N_NET256_XI39/MM2437_g N_VSS_XI39/MM2437_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2518 N_NET416_XI39/MM2518_d N_NET387_XI39/MM2518_g N_VSS_XI39/MM2518_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2501 XI39/NET11442 N_NET388_XI39/MM2501_g N_VSS_XI39/MM2501_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2537 N_NET416_XI39/MM2537_d N_NET389_XI39/MM2537_g N_VSS_XI39/MM2537_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2548 XI39/NET11630 N_NET390_XI39/MM2548_g N_VSS_XI39/MM2548_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2217 N_NET416_XI39/MM2217_d N_NET391_XI39/MM2217_g N_VSS_XI39/MM2217_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2228 XI39/NET10442 N_NET262_XI39/MM2228_g N_VSS_XI39/MM2228_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2198 N_NET416_XI39/MM2198_d N_NET263_XI39/MM2198_g N_VSS_XI39/MM2198_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2181 XI39/NET10622 N_NET264_XI39/MM2181_g N_VSS_XI39/MM2181_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2262 N_NET416_XI39/MM2262_d N_NET265_XI39/MM2262_g N_VSS_XI39/MM2262_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2245 XI39/NET10374 N_NET396_XI39/MM2245_g N_VSS_XI39/MM2245_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2281 N_NET416_XI39/MM2281_d N_NET267_XI39/MM2281_g N_VSS_XI39/MM2281_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2292 XI39/NET10194 N_NET268_XI39/MM2292_g N_VSS_XI39/MM2292_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2134 N_NET416_XI39/MM2134_d N_NET269_XI39/MM2134_g N_VSS_XI39/MM2134_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2117 XI39/NET9858 N_NET270_XI39/MM2117_g N_VSS_XI39/MM2117_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2153 N_NET416_XI39/MM2153_d N_NET401_XI39/MM2153_g N_VSS_XI39/MM2153_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2164 XI39/NET9678 N_NET272_XI39/MM2164_g N_VSS_XI39/MM2164_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2089 N_NET416_XI39/MM2089_d N_NET273_XI39/MM2089_g N_VSS_XI39/MM2089_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2100 XI39/NET9930 N_NET404_XI39/MM2100_g N_VSS_XI39/MM2100_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2070 N_NET416_XI39/MM2070_d N_NET405_XI39/MM2070_g N_VSS_XI39/MM2070_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4 XI39/NET10058 N_NET0390_XI39/MM4_g N_VSS_XI39/MM4_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI54/XI1/XI6/MM1 N_XI54/XI1/NET2_XI54/XI1/XI6/MM1_d N_NET061_XI54/XI1/XI6/MM1_g
+ N_VSS_XI54/XI1/XI6/MM1_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI39/MM3418 XI39/NET5550 N_NET0133_XI39/MM3418_g N_VSS_XI39/MM3418_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3400 N_NET417_XI39/MM3400_d N_NET280_XI39/MM3400_g N_VSS_XI39/MM3400_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3431 XI39/NET5498 N_NET281_XI39/MM3431_g N_VSS_XI39/MM3431_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3446 N_NET417_XI39/MM3446_d N_NET282_XI39/MM3446_g N_VSS_XI39/MM3446_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3368 XI39/NET5750 N_NET153_XI39/MM3368_g N_VSS_XI39/MM3368_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3383 N_NET417_XI39/MM3383_d N_NET284_XI39/MM3383_g N_VSS_XI39/MM3383_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3353 XI39/NET3510 N_NET285_XI39/MM3353_g N_VSS_XI39/MM3353_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3336 N_NET417_XI39/MM3336_d N_NET286_XI39/MM3336_g N_VSS_XI39/MM3336_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3495 XI39/NET5242 N_NET287_XI39/MM3495_g N_VSS_XI39/MM3495_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3510 N_NET417_XI39/MM3510_d N_NET158_XI39/MM3510_g N_VSS_XI39/MM3510_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3480 XI39/NET5302 N_NET159_XI39/MM3480_g N_VSS_XI39/MM3480_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3463 N_NET417_XI39/MM3463_d N_NET160_XI39/MM3463_g N_VSS_XI39/MM3463_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3544 XI39/NET5046 N_NET291_XI39/MM3544_g N_VSS_XI39/MM3544_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3527 N_NET417_XI39/MM3527_d N_NET162_XI39/MM3527_g N_VSS_XI39/MM3527_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3559 XI39/NET4986 N_NET293_XI39/MM3559_g N_VSS_XI39/MM3559_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3574 N_NET417_XI39/MM3574_d N_NET294_XI39/MM3574_g N_VSS_XI39/MM3574_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3240 XI39/NET3962 N_NET295_XI39/MM3240_g N_VSS_XI39/MM3240_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3255 N_NET417_XI39/MM3255_d N_NET296_XI39/MM3255_g N_VSS_XI39/MM3255_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3225 XI39/NET4022 N_NET297_XI39/MM3225_g N_VSS_XI39/MM3225_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3208 N_NET417_XI39/MM3208_d N_NET298_XI39/MM3208_g N_VSS_XI39/MM3208_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3289 XI39/NET3766 N_NET299_XI39/MM3289_g N_VSS_XI39/MM3289_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3272 N_NET417_XI39/MM3272_d N_NET170_XI39/MM3272_g N_VSS_XI39/MM3272_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3304 XI39/NET3706 N_NET171_XI39/MM3304_g N_VSS_XI39/MM3304_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3319 N_NET417_XI39/MM3319_d N_NET172_XI39/MM3319_g N_VSS_XI39/MM3319_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3161 XI39/NET4278 N_NET303_XI39/MM3161_g N_VSS_XI39/MM3161_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3144 N_NET417_XI39/MM3144_d N_NET304_XI39/MM3144_g N_VSS_XI39/MM3144_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3176 XI39/NET4218 N_NET305_XI39/MM3176_g N_VSS_XI39/MM3176_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3191 N_NET417_XI39/MM3191_d N_NET306_XI39/MM3191_g N_VSS_XI39/MM3191_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3112 XI39/NET4474 N_NET307_XI39/MM3112_g N_VSS_XI39/MM3112_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3127 N_NET417_XI39/MM3127_d N_NET308_XI39/MM3127_g N_VSS_XI39/MM3127_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3097 XI39/NET4534 N_NET309_XI39/MM3097_g N_VSS_XI39/MM3097_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3080 N_NET417_XI39/MM3080_d N_NET310_XI39/MM3080_g N_VSS_XI39/MM3080_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3841 XI39/NET6158 N_NET311_XI39/MM3841_g N_VSS_XI39/MM3841_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3856 N_NET417_XI39/MM3856_d N_NET312_XI39/MM3856_g N_VSS_XI39/MM3856_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3988 XI39/NET7366 N_NET313_XI39/MM3988_g N_VSS_XI39/MM3988_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3971 N_NET417_XI39/MM3971_d N_NET314_XI39/MM3971_g N_VSS_XI39/MM3971_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3890 XI39/NET5962 N_NET315_XI39/MM3890_g N_VSS_XI39/MM3890_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3873 N_NET417_XI39/MM3873_d N_NET316_XI39/MM3873_g N_VSS_XI39/MM3873_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3905 XI39/NET5902 N_NET317_XI39/MM3905_g N_VSS_XI39/MM3905_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3920 N_NET417_XI39/MM3920_d N_NET318_XI39/MM3920_g N_VSS_XI39/MM3920_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4068 XI39/NET7046 N_NET319_XI39/MM4068_g N_VSS_XI39/MM4068_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4051 N_NET417_XI39/MM4051_d N_NET320_XI39/MM4051_g N_VSS_XI39/MM4051_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3943 XI39/NET7546 N_NET321_XI39/MM3943_g N_VSS_XI39/MM3943_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3954 N_NET417_XI39/MM3954_d N_NET192_XI39/MM3954_g N_VSS_XI39/MM3954_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4019 XI39/NET7242 N_NET193_XI39/MM4019_g N_VSS_XI39/MM4019_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4034 N_NET417_XI39/MM4034_d N_NET194_XI39/MM4034_g N_VSS_XI39/MM4034_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4010 XI39/NET7278 N_NET195_XI39/MM4010_g N_VSS_XI39/MM4010_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4081 N_NET417_XI39/MM4081_d N_NET196_XI39/MM4081_g N_VSS_XI39/MM4081_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3800 XI39/NET6322 N_NET197_XI39/MM3800_g N_VSS_XI39/MM3800_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3783 N_NET417_XI39/MM3783_d N_NET198_XI39/MM3783_g N_VSS_XI39/MM3783_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3815 XI39/NET6262 N_NET199_XI39/MM3815_g N_VSS_XI39/MM3815_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3830 N_NET417_XI39/MM3830_d N_NET200_XI39/MM3830_g N_VSS_XI39/MM3830_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3751 XI39/NET6518 N_NET331_XI39/MM3751_g N_VSS_XI39/MM3751_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3766 N_NET417_XI39/MM3766_d N_NET332_XI39/MM3766_g N_VSS_XI39/MM3766_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3736 XI39/NET6578 N_NET203_XI39/MM3736_g N_VSS_XI39/MM3736_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3719 N_NET417_XI39/MM3719_d N_NET204_XI39/MM3719_g N_VSS_XI39/MM3719_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3623 XI39/NET4730 N_NET205_XI39/MM3623_g N_VSS_XI39/MM3623_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3638 N_NET417_XI39/MM3638_d N_NET206_XI39/MM3638_g N_VSS_XI39/MM3638_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3608 XI39/NET4790 N_NET207_XI39/MM3608_g N_VSS_XI39/MM3608_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3591 N_NET417_XI39/MM3591_d N_NET338_XI39/MM3591_g N_VSS_XI39/MM3591_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3672 XI39/NET6834 N_NET339_XI39/MM3672_g N_VSS_XI39/MM3672_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3655 N_NET417_XI39/MM3655_d N_NET340_XI39/MM3655_g N_VSS_XI39/MM3655_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3704 XI39/NET6706 N_NET211_XI39/MM3704_g N_VSS_XI39/MM3704_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3695 N_NET417_XI39/MM3695_d N_NET212_XI39/MM3695_g N_VSS_XI39/MM3695_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2728 XI39/NET8950 N_NET214_XI39/MM2728_g N_VSS_XI39/MM2728_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2743 N_NET417_XI39/MM2743_d N_NET215_XI39/MM2743_g N_VSS_XI39/MM2743_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2713 XI39/NET9010 N_NET216_XI39/MM2713_g N_VSS_XI39/MM2713_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2696 N_NET417_XI39/MM2696_d N_NET346_XI39/MM2696_g N_VSS_XI39/MM2696_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2777 XI39/NET8758 N_NET347_XI39/MM2777_g N_VSS_XI39/MM2777_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2760 N_NET417_XI39/MM2760_d N_NET348_XI39/MM2760_g N_VSS_XI39/MM2760_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2792 XI39/NET8698 N_NET349_XI39/MM2792_g N_VSS_XI39/MM2792_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2807 N_NET417_XI39/MM2807_d N_NET350_XI39/MM2807_g N_VSS_XI39/MM2807_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2649 XI39/NET9266 N_NET351_XI39/MM2649_g N_VSS_XI39/MM2649_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2632 N_NET417_XI39/MM2632_d N_NET352_XI39/MM2632_g N_VSS_XI39/MM2632_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2664 XI39/NET9206 N_NET224_XI39/MM2664_g N_VSS_XI39/MM2664_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2679 N_NET417_XI39/MM2679_d N_NET225_XI39/MM2679_g N_VSS_XI39/MM2679_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2600 XI39/NET9462 N_NET226_XI39/MM2600_g N_VSS_XI39/MM2600_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2615 N_NET417_XI39/MM2615_d N_NET356_XI39/MM2615_g N_VSS_XI39/MM2615_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2585 XI39/NET9522 N_NET357_XI39/MM2585_g N_VSS_XI39/MM2585_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2568 N_NET417_XI39/MM2568_d N_NET358_XI39/MM2568_g N_VSS_XI39/MM2568_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2905 XI39/NET8246 N_NET230_XI39/MM2905_g N_VSS_XI39/MM2905_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2888 N_NET417_XI39/MM2888_d N_NET360_XI39/MM2888_g N_VSS_XI39/MM2888_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2920 XI39/NET8186 N_NET361_XI39/MM2920_g N_VSS_XI39/MM2920_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2935 N_NET417_XI39/MM2935_d N_NET233_XI39/MM2935_g N_VSS_XI39/MM2935_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2856 XI39/NET8442 N_NET234_XI39/MM2856_g N_VSS_XI39/MM2856_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2871 N_NET417_XI39/MM2871_d N_NET235_XI39/MM2871_g N_VSS_XI39/MM2871_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2841 XI39/NET8502 N_NET365_XI39/MM2841_g N_VSS_XI39/MM2841_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2824 N_NET417_XI39/MM2824_d N_NET366_XI39/MM2824_g N_VSS_XI39/MM2824_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2984 XI39/NET7930 N_NET367_XI39/MM2984_g N_VSS_XI39/MM2984_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2999 N_NET417_XI39/MM2999_d N_NET368_XI39/MM2999_g N_VSS_XI39/MM2999_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2969 XI39/NET7990 N_NET369_XI39/MM2969_g N_VSS_XI39/MM2969_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2952 N_NET417_XI39/MM2952_d N_NET370_XI39/MM2952_g N_VSS_XI39/MM2952_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3033 XI39/NET7734 N_NET371_XI39/MM3033_g N_VSS_XI39/MM3033_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3016 N_NET417_XI39/MM3016_d N_NET242_XI39/MM3016_g N_VSS_XI39/MM3016_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3048 XI39/NET7674 N_NET373_XI39/MM3048_g N_VSS_XI39/MM3048_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3063 N_NET417_XI39/MM3063_d N_NET244_XI39/MM3063_g N_VSS_XI39/MM3063_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2387 XI39/NET10674 N_NET375_XI39/MM2387_g N_VSS_XI39/MM2387_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2376 N_NET417_XI39/MM2376_d N_NET376_XI39/MM2376_g N_VSS_XI39/MM2376_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2408 XI39/NET11238 N_NET377_XI39/MM2408_g N_VSS_XI39/MM2408_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2423 N_NET417_XI39/MM2423_d N_NET378_XI39/MM2423_g N_VSS_XI39/MM2423_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2344 XI39/NET10846 N_NET379_XI39/MM2344_g N_VSS_XI39/MM2344_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2359 N_NET417_XI39/MM2359_d N_NET380_XI39/MM2359_g N_VSS_XI39/MM2359_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2329 XI39/NET10906 N_NET381_XI39/MM2329_g N_VSS_XI39/MM2329_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2312 N_NET417_XI39/MM2312_d N_NET382_XI39/MM2312_g N_VSS_XI39/MM2312_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2474 XI39/NET11550 N_NET383_XI39/MM2474_g N_VSS_XI39/MM2474_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2487 N_NET417_XI39/MM2487_d N_NET384_XI39/MM2487_g N_VSS_XI39/MM2487_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2457 XI39/NET11042 N_NET385_XI39/MM2457_g N_VSS_XI39/MM2457_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2440 N_NET417_XI39/MM2440_d N_NET256_XI39/MM2440_g N_VSS_XI39/MM2440_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2521 XI39/NET11362 N_NET387_XI39/MM2521_g N_VSS_XI39/MM2521_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2504 N_NET417_XI39/MM2504_d N_NET388_XI39/MM2504_g N_VSS_XI39/MM2504_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2530 XI39/NET11326 N_NET389_XI39/MM2530_g N_VSS_XI39/MM2530_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2551 N_NET417_XI39/MM2551_d N_NET390_XI39/MM2551_g N_VSS_XI39/MM2551_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2216 XI39/NET10486 N_NET391_XI39/MM2216_g N_VSS_XI39/MM2216_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2231 N_NET417_XI39/MM2231_d N_NET262_XI39/MM2231_g N_VSS_XI39/MM2231_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2201 XI39/NET10546 N_NET263_XI39/MM2201_g N_VSS_XI39/MM2201_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2184 N_NET417_XI39/MM2184_d N_NET264_XI39/MM2184_g N_VSS_XI39/MM2184_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2265 XI39/NET10298 N_NET265_XI39/MM2265_g N_VSS_XI39/MM2265_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2248 N_NET417_XI39/MM2248_d N_NET396_XI39/MM2248_g N_VSS_XI39/MM2248_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2280 XI39/NET10238 N_NET267_XI39/MM2280_g N_VSS_XI39/MM2280_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2295 N_NET417_XI39/MM2295_d N_NET268_XI39/MM2295_g N_VSS_XI39/MM2295_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2139 XI39/NET9774 N_NET269_XI39/MM2139_g N_VSS_XI39/MM2139_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2120 N_NET417_XI39/MM2120_d N_NET270_XI39/MM2120_g N_VSS_XI39/MM2120_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2152 XI39/NET9722 N_NET401_XI39/MM2152_g N_VSS_XI39/MM2152_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2167 N_NET417_XI39/MM2167_d N_NET272_XI39/MM2167_g N_VSS_XI39/MM2167_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2088 XI39/NET9974 N_NET273_XI39/MM2088_g N_VSS_XI39/MM2088_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2103 N_NET417_XI39/MM2103_d N_NET404_XI39/MM2103_g N_VSS_XI39/MM2103_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2071 XI39/NET10034 N_NET405_XI39/MM2071_g N_VSS_XI39/MM2071_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM7 N_NET417_XI39/MM7_d N_NET0390_XI39/MM7_g N_VSS_XI39/MM7_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI29/XI1/MM39 N_NET481_XI29/XI1/MM39_d N_XI29/XI1/NET195_XI29/XI1/MM39_g
+ N_NET065_XI29/XI1/MM39_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI29/XI1/XI8/MM1 N_XI29/XI1/NET195_XI29/XI1/XI8/MM1_d
+ N_NET470_XI29/XI1/XI8/MM1_g N_VSS_XI29/XI1/XI8/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI29/XI1/MM40 N_NET482_XI29/XI1/MM40_d N_XI29/XI1/NET199_XI29/XI1/MM40_g
+ N_NET065_XI29/XI1/MM40_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI29/XI1/XI9/MM1 N_XI29/XI1/NET199_XI29/XI1/XI9/MM1_d
+ N_NET469_XI29/XI1/XI9/MM1_g N_VSS_XI29/XI1/XI9/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI39/MM3415 N_NET481_XI39/MM3415_d N_NET0133_XI39/MM3415_g N_VSS_XI39/MM3415_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3399 XI39/NET5626 N_NET280_XI39/MM3399_g N_VSS_XI39/MM3399_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3430 N_NET481_XI39/MM3430_d N_NET281_XI39/MM3430_g N_VSS_XI39/MM3430_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3445 XI39/NET5442 N_NET282_XI39/MM3445_g N_VSS_XI39/MM3445_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3367 N_NET481_XI39/MM3367_d N_NET153_XI39/MM3367_g N_VSS_XI39/MM3367_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3382 XI39/NET5694 N_NET284_XI39/MM3382_g N_VSS_XI39/MM3382_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3352 N_NET481_XI39/MM3352_d N_NET285_XI39/MM3352_g N_VSS_XI39/MM3352_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3343 XI39/NET3550 N_NET286_XI39/MM3343_g N_VSS_XI39/MM3343_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3494 N_NET481_XI39/MM3494_d N_NET287_XI39/MM3494_g N_VSS_XI39/MM3494_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3509 XI39/NET5186 N_NET158_XI39/MM3509_g N_VSS_XI39/MM3509_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3479 N_NET481_XI39/MM3479_d N_NET159_XI39/MM3479_g N_VSS_XI39/MM3479_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3462 XI39/NET5374 N_NET160_XI39/MM3462_g N_VSS_XI39/MM3462_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3543 N_NET481_XI39/MM3543_d N_NET291_XI39/MM3543_g N_VSS_XI39/MM3543_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3526 XI39/NET5118 N_NET162_XI39/MM3526_g N_VSS_XI39/MM3526_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3558 N_NET481_XI39/MM3558_d N_NET293_XI39/MM3558_g N_VSS_XI39/MM3558_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3573 XI39/NET4930 N_NET294_XI39/MM3573_g N_VSS_XI39/MM3573_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3239 N_NET481_XI39/MM3239_d N_NET295_XI39/MM3239_g N_VSS_XI39/MM3239_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3254 XI39/NET3906 N_NET296_XI39/MM3254_g N_VSS_XI39/MM3254_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3224 N_NET481_XI39/MM3224_d N_NET297_XI39/MM3224_g N_VSS_XI39/MM3224_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3207 XI39/NET4094 N_NET298_XI39/MM3207_g N_VSS_XI39/MM3207_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3288 N_NET481_XI39/MM3288_d N_NET299_XI39/MM3288_g N_VSS_XI39/MM3288_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3271 XI39/NET3838 N_NET170_XI39/MM3271_g N_VSS_XI39/MM3271_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3303 N_NET481_XI39/MM3303_d N_NET171_XI39/MM3303_g N_VSS_XI39/MM3303_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3318 XI39/NET3650 N_NET172_XI39/MM3318_g N_VSS_XI39/MM3318_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3160 N_NET481_XI39/MM3160_d N_NET303_XI39/MM3160_g N_VSS_XI39/MM3160_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3143 XI39/NET4350 N_NET304_XI39/MM3143_g N_VSS_XI39/MM3143_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3175 N_NET481_XI39/MM3175_d N_NET305_XI39/MM3175_g N_VSS_XI39/MM3175_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3190 XI39/NET4162 N_NET306_XI39/MM3190_g N_VSS_XI39/MM3190_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3111 N_NET481_XI39/MM3111_d N_NET307_XI39/MM3111_g N_VSS_XI39/MM3111_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3126 XI39/NET4418 N_NET308_XI39/MM3126_g N_VSS_XI39/MM3126_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3096 N_NET481_XI39/MM3096_d N_NET309_XI39/MM3096_g N_VSS_XI39/MM3096_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3079 XI39/NET4606 N_NET310_XI39/MM3079_g N_VSS_XI39/MM3079_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3840 N_NET481_XI39/MM3840_d N_NET311_XI39/MM3840_g N_VSS_XI39/MM3840_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3855 XI39/NET6102 N_NET312_XI39/MM3855_g N_VSS_XI39/MM3855_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3987 N_NET481_XI39/MM3987_d N_NET313_XI39/MM3987_g N_VSS_XI39/MM3987_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3970 XI39/NET7438 N_NET314_XI39/MM3970_g N_VSS_XI39/MM3970_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3889 N_NET481_XI39/MM3889_d N_NET315_XI39/MM3889_g N_VSS_XI39/MM3889_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3872 XI39/NET6034 N_NET316_XI39/MM3872_g N_VSS_XI39/MM3872_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3904 N_NET481_XI39/MM3904_d N_NET317_XI39/MM3904_g N_VSS_XI39/MM3904_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3919 XI39/NET5846 N_NET318_XI39/MM3919_g N_VSS_XI39/MM3919_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4067 N_NET481_XI39/MM4067_d N_NET319_XI39/MM4067_g N_VSS_XI39/MM4067_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4050 XI39/NET7118 N_NET320_XI39/MM4050_g N_VSS_XI39/MM4050_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3938 N_NET481_XI39/MM3938_d N_NET321_XI39/MM3938_g N_VSS_XI39/MM3938_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3953 XI39/NET7506 N_NET192_XI39/MM3953_g N_VSS_XI39/MM3953_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4018 N_NET481_XI39/MM4018_d N_NET193_XI39/MM4018_g N_VSS_XI39/MM4018_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4033 XI39/NET7186 N_NET194_XI39/MM4033_g N_VSS_XI39/MM4033_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4003 N_NET481_XI39/MM4003_d N_NET195_XI39/MM4003_g N_VSS_XI39/MM4003_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4080 XI39/NET6998 N_NET196_XI39/MM4080_g N_VSS_XI39/MM4080_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3799 N_NET481_XI39/MM3799_d N_NET197_XI39/MM3799_g N_VSS_XI39/MM3799_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3782 XI39/NET6394 N_NET198_XI39/MM3782_g N_VSS_XI39/MM3782_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3814 N_NET481_XI39/MM3814_d N_NET199_XI39/MM3814_g N_VSS_XI39/MM3814_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3829 XI39/NET6206 N_NET200_XI39/MM3829_g N_VSS_XI39/MM3829_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3750 N_NET481_XI39/MM3750_d N_NET331_XI39/MM3750_g N_VSS_XI39/MM3750_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3765 XI39/NET6462 N_NET332_XI39/MM3765_g N_VSS_XI39/MM3765_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3735 N_NET481_XI39/MM3735_d N_NET203_XI39/MM3735_g N_VSS_XI39/MM3735_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3718 XI39/NET6650 N_NET204_XI39/MM3718_g N_VSS_XI39/MM3718_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3622 N_NET481_XI39/MM3622_d N_NET205_XI39/MM3622_g N_VSS_XI39/MM3622_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3637 XI39/NET4674 N_NET206_XI39/MM3637_g N_VSS_XI39/MM3637_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3607 N_NET481_XI39/MM3607_d N_NET207_XI39/MM3607_g N_VSS_XI39/MM3607_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3590 XI39/NET4862 N_NET338_XI39/MM3590_g N_VSS_XI39/MM3590_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3671 N_NET481_XI39/MM3671_d N_NET339_XI39/MM3671_g N_VSS_XI39/MM3671_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3654 XI39/NET6906 N_NET340_XI39/MM3654_g N_VSS_XI39/MM3654_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3687 N_NET481_XI39/MM3687_d N_NET211_XI39/MM3687_g N_VSS_XI39/MM3687_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3694 XI39/NET6746 N_NET212_XI39/MM3694_g N_VSS_XI39/MM3694_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2727 N_NET481_XI39/MM2727_d N_NET214_XI39/MM2727_g N_VSS_XI39/MM2727_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2742 XI39/NET8898 N_NET215_XI39/MM2742_g N_VSS_XI39/MM2742_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2712 N_NET481_XI39/MM2712_d N_NET216_XI39/MM2712_g N_VSS_XI39/MM2712_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2695 XI39/NET9082 N_NET346_XI39/MM2695_g N_VSS_XI39/MM2695_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2776 N_NET481_XI39/MM2776_d N_NET347_XI39/MM2776_g N_VSS_XI39/MM2776_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2759 XI39/NET8830 N_NET348_XI39/MM2759_g N_VSS_XI39/MM2759_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2791 N_NET481_XI39/MM2791_d N_NET349_XI39/MM2791_g N_VSS_XI39/MM2791_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2806 XI39/NET8642 N_NET350_XI39/MM2806_g N_VSS_XI39/MM2806_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2648 N_NET481_XI39/MM2648_d N_NET351_XI39/MM2648_g N_VSS_XI39/MM2648_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2631 XI39/NET9338 N_NET352_XI39/MM2631_g N_VSS_XI39/MM2631_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2663 N_NET481_XI39/MM2663_d N_NET224_XI39/MM2663_g N_VSS_XI39/MM2663_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2678 XI39/NET9150 N_NET225_XI39/MM2678_g N_VSS_XI39/MM2678_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2599 N_NET481_XI39/MM2599_d N_NET226_XI39/MM2599_g N_VSS_XI39/MM2599_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2614 XI39/NET9406 N_NET356_XI39/MM2614_g N_VSS_XI39/MM2614_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2584 N_NET481_XI39/MM2584_d N_NET357_XI39/MM2584_g N_VSS_XI39/MM2584_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2567 XI39/NET9594 N_NET358_XI39/MM2567_g N_VSS_XI39/MM2567_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2904 N_NET481_XI39/MM2904_d N_NET230_XI39/MM2904_g N_VSS_XI39/MM2904_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2887 XI39/NET8318 N_NET360_XI39/MM2887_g N_VSS_XI39/MM2887_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2919 N_NET481_XI39/MM2919_d N_NET361_XI39/MM2919_g N_VSS_XI39/MM2919_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2934 XI39/NET8130 N_NET233_XI39/MM2934_g N_VSS_XI39/MM2934_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2855 N_NET481_XI39/MM2855_d N_NET234_XI39/MM2855_g N_VSS_XI39/MM2855_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2870 XI39/NET8386 N_NET235_XI39/MM2870_g N_VSS_XI39/MM2870_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2840 N_NET481_XI39/MM2840_d N_NET365_XI39/MM2840_g N_VSS_XI39/MM2840_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2823 XI39/NET8574 N_NET366_XI39/MM2823_g N_VSS_XI39/MM2823_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2983 N_NET481_XI39/MM2983_d N_NET367_XI39/MM2983_g N_VSS_XI39/MM2983_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2998 XI39/NET7874 N_NET368_XI39/MM2998_g N_VSS_XI39/MM2998_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2968 N_NET481_XI39/MM2968_d N_NET369_XI39/MM2968_g N_VSS_XI39/MM2968_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2951 XI39/NET8062 N_NET370_XI39/MM2951_g N_VSS_XI39/MM2951_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3032 N_NET481_XI39/MM3032_d N_NET371_XI39/MM3032_g N_VSS_XI39/MM3032_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3015 XI39/NET7806 N_NET242_XI39/MM3015_g N_VSS_XI39/MM3015_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3047 N_NET481_XI39/MM3047_d N_NET373_XI39/MM3047_g N_VSS_XI39/MM3047_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3062 XI39/NET7618 N_NET244_XI39/MM3062_g N_VSS_XI39/MM3062_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2392 N_NET481_XI39/MM2392_d N_NET375_XI39/MM2392_g N_VSS_XI39/MM2392_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2375 XI39/NET10722 N_NET376_XI39/MM2375_g N_VSS_XI39/MM2375_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2407 N_NET481_XI39/MM2407_d N_NET377_XI39/MM2407_g N_VSS_XI39/MM2407_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2422 XI39/NET11182 N_NET378_XI39/MM2422_g N_VSS_XI39/MM2422_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2343 N_NET481_XI39/MM2343_d N_NET379_XI39/MM2343_g N_VSS_XI39/MM2343_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2358 XI39/NET10790 N_NET380_XI39/MM2358_g N_VSS_XI39/MM2358_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2328 N_NET481_XI39/MM2328_d N_NET381_XI39/MM2328_g N_VSS_XI39/MM2328_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2311 XI39/NET10978 N_NET382_XI39/MM2311_g N_VSS_XI39/MM2311_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2471 N_NET481_XI39/MM2471_d N_NET383_XI39/MM2471_g N_VSS_XI39/MM2471_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2486 XI39/NET11502 N_NET384_XI39/MM2486_g N_VSS_XI39/MM2486_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2456 N_NET481_XI39/MM2456_d N_NET385_XI39/MM2456_g N_VSS_XI39/MM2456_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2439 XI39/NET11114 N_NET256_XI39/MM2439_g N_VSS_XI39/MM2439_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2520 N_NET481_XI39/MM2520_d N_NET387_XI39/MM2520_g N_VSS_XI39/MM2520_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2503 XI39/NET11434 N_NET388_XI39/MM2503_g N_VSS_XI39/MM2503_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2535 N_NET481_XI39/MM2535_d N_NET389_XI39/MM2535_g N_VSS_XI39/MM2535_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2550 XI39/NET11622 N_NET390_XI39/MM2550_g N_VSS_XI39/MM2550_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2215 N_NET481_XI39/MM2215_d N_NET391_XI39/MM2215_g N_VSS_XI39/MM2215_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2230 XI39/NET10434 N_NET262_XI39/MM2230_g N_VSS_XI39/MM2230_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2200 N_NET481_XI39/MM2200_d N_NET263_XI39/MM2200_g N_VSS_XI39/MM2200_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2183 XI39/NET10614 N_NET264_XI39/MM2183_g N_VSS_XI39/MM2183_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2264 N_NET481_XI39/MM2264_d N_NET265_XI39/MM2264_g N_VSS_XI39/MM2264_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2247 XI39/NET10366 N_NET396_XI39/MM2247_g N_VSS_XI39/MM2247_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2279 N_NET481_XI39/MM2279_d N_NET267_XI39/MM2279_g N_VSS_XI39/MM2279_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2294 XI39/NET10186 N_NET268_XI39/MM2294_g N_VSS_XI39/MM2294_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2136 N_NET481_XI39/MM2136_d N_NET269_XI39/MM2136_g N_VSS_XI39/MM2136_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2119 XI39/NET9850 N_NET270_XI39/MM2119_g N_VSS_XI39/MM2119_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2151 N_NET481_XI39/MM2151_d N_NET401_XI39/MM2151_g N_VSS_XI39/MM2151_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2166 XI39/NET9670 N_NET272_XI39/MM2166_g N_VSS_XI39/MM2166_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2087 N_NET481_XI39/MM2087_d N_NET273_XI39/MM2087_g N_VSS_XI39/MM2087_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2102 XI39/NET9922 N_NET404_XI39/MM2102_g N_VSS_XI39/MM2102_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2072 N_NET481_XI39/MM2072_d N_NET405_XI39/MM2072_g N_VSS_XI39/MM2072_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM10 XI39/NET10082 N_NET0390_XI39/MM10_g N_VSS_XI39/MM10_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI54/XI1/XI8/XI3/MM3 N_XI54/XI1/XI8/XI3/NET13_XI54/XI1/XI8/XI3/MM3_d
+ N_XI54/XI1/NET2_XI54/XI1/XI8/XI3/MM3_g N_VSS_XI54/XI1/XI8/XI3/MM3_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=1.68025e-13
+ AS=2.303e-13 PD=7.15e-07 PS=1.45e-06
mXI54/XI1/XI7/XI3/MM3 N_XI54/XI1/XI7/XI3/NET13_XI54/XI1/XI7/XI3/MM3_d
+ N_NET061_XI54/XI1/XI7/XI3/MM3_g N_VSS_XI54/XI1/XI7/XI3/MM3_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=1.68025e-13
+ AS=2.303e-13 PD=7.15e-07 PS=1.45e-06
mXI39/MM3412 XI39/NET5574 N_NET0133_XI39/MM3412_g N_VSS_XI39/MM3412_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3398 N_NET482_XI39/MM3398_d N_NET280_XI39/MM3398_g N_VSS_XI39/MM3398_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3433 XI39/NET5490 N_NET281_XI39/MM3433_g N_VSS_XI39/MM3433_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3448 N_NET482_XI39/MM3448_d N_NET282_XI39/MM3448_g N_VSS_XI39/MM3448_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3370 XI39/NET5742 N_NET153_XI39/MM3370_g N_VSS_XI39/MM3370_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3385 N_NET482_XI39/MM3385_d N_NET284_XI39/MM3385_g N_VSS_XI39/MM3385_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3355 XI39/NET3502 N_NET285_XI39/MM3355_g N_VSS_XI39/MM3355_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3334 N_NET482_XI39/MM3334_d N_NET286_XI39/MM3334_g N_VSS_XI39/MM3334_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3497 XI39/NET5234 N_NET287_XI39/MM3497_g N_VSS_XI39/MM3497_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3512 N_NET482_XI39/MM3512_d N_NET158_XI39/MM3512_g N_VSS_XI39/MM3512_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3482 XI39/NET5294 N_NET159_XI39/MM3482_g N_VSS_XI39/MM3482_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3461 N_NET482_XI39/MM3461_d N_NET160_XI39/MM3461_g N_VSS_XI39/MM3461_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3546 XI39/NET5038 N_NET291_XI39/MM3546_g N_VSS_XI39/MM3546_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3525 N_NET482_XI39/MM3525_d N_NET162_XI39/MM3525_g N_VSS_XI39/MM3525_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3561 XI39/NET4978 N_NET293_XI39/MM3561_g N_VSS_XI39/MM3561_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3576 N_NET482_XI39/MM3576_d N_NET294_XI39/MM3576_g N_VSS_XI39/MM3576_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3242 XI39/NET3954 N_NET295_XI39/MM3242_g N_VSS_XI39/MM3242_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3257 N_NET482_XI39/MM3257_d N_NET296_XI39/MM3257_g N_VSS_XI39/MM3257_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3227 XI39/NET4014 N_NET297_XI39/MM3227_g N_VSS_XI39/MM3227_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3206 N_NET482_XI39/MM3206_d N_NET298_XI39/MM3206_g N_VSS_XI39/MM3206_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3291 XI39/NET3758 N_NET299_XI39/MM3291_g N_VSS_XI39/MM3291_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3270 N_NET482_XI39/MM3270_d N_NET170_XI39/MM3270_g N_VSS_XI39/MM3270_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3306 XI39/NET3698 N_NET171_XI39/MM3306_g N_VSS_XI39/MM3306_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3321 N_NET482_XI39/MM3321_d N_NET172_XI39/MM3321_g N_VSS_XI39/MM3321_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3163 XI39/NET4270 N_NET303_XI39/MM3163_g N_VSS_XI39/MM3163_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3142 N_NET482_XI39/MM3142_d N_NET304_XI39/MM3142_g N_VSS_XI39/MM3142_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3178 XI39/NET4210 N_NET305_XI39/MM3178_g N_VSS_XI39/MM3178_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3193 N_NET482_XI39/MM3193_d N_NET306_XI39/MM3193_g N_VSS_XI39/MM3193_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3114 XI39/NET4466 N_NET307_XI39/MM3114_g N_VSS_XI39/MM3114_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3129 N_NET482_XI39/MM3129_d N_NET308_XI39/MM3129_g N_VSS_XI39/MM3129_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3099 XI39/NET4526 N_NET309_XI39/MM3099_g N_VSS_XI39/MM3099_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3078 N_NET482_XI39/MM3078_d N_NET310_XI39/MM3078_g N_VSS_XI39/MM3078_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3843 XI39/NET6150 N_NET311_XI39/MM3843_g N_VSS_XI39/MM3843_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3858 N_NET482_XI39/MM3858_d N_NET312_XI39/MM3858_g N_VSS_XI39/MM3858_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3990 XI39/NET7358 N_NET313_XI39/MM3990_g N_VSS_XI39/MM3990_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3969 N_NET482_XI39/MM3969_d N_NET314_XI39/MM3969_g N_VSS_XI39/MM3969_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3892 XI39/NET5954 N_NET315_XI39/MM3892_g N_VSS_XI39/MM3892_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3871 N_NET482_XI39/MM3871_d N_NET316_XI39/MM3871_g N_VSS_XI39/MM3871_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3907 XI39/NET5894 N_NET317_XI39/MM3907_g N_VSS_XI39/MM3907_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3922 N_NET482_XI39/MM3922_d N_NET318_XI39/MM3922_g N_VSS_XI39/MM3922_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4070 XI39/NET7038 N_NET319_XI39/MM4070_g N_VSS_XI39/MM4070_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4049 N_NET482_XI39/MM4049_d N_NET320_XI39/MM4049_g N_VSS_XI39/MM4049_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3945 XI39/NET7538 N_NET321_XI39/MM3945_g N_VSS_XI39/MM3945_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3956 N_NET482_XI39/MM3956_d N_NET192_XI39/MM3956_g N_VSS_XI39/MM3956_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4021 XI39/NET7234 N_NET193_XI39/MM4021_g N_VSS_XI39/MM4021_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4036 N_NET482_XI39/MM4036_d N_NET194_XI39/MM4036_g N_VSS_XI39/MM4036_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4090 XI39/NET6958 N_NET195_XI39/MM4090_g N_VSS_XI39/MM4090_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4079 N_NET482_XI39/MM4079_d N_NET196_XI39/MM4079_g N_VSS_XI39/MM4079_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3802 XI39/NET6314 N_NET197_XI39/MM3802_g N_VSS_XI39/MM3802_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3781 N_NET482_XI39/MM3781_d N_NET198_XI39/MM3781_g N_VSS_XI39/MM3781_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3817 XI39/NET6254 N_NET199_XI39/MM3817_g N_VSS_XI39/MM3817_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3832 N_NET482_XI39/MM3832_d N_NET200_XI39/MM3832_g N_VSS_XI39/MM3832_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3753 XI39/NET6510 N_NET331_XI39/MM3753_g N_VSS_XI39/MM3753_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3768 N_NET482_XI39/MM3768_d N_NET332_XI39/MM3768_g N_VSS_XI39/MM3768_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3738 XI39/NET6570 N_NET203_XI39/MM3738_g N_VSS_XI39/MM3738_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3717 N_NET482_XI39/MM3717_d N_NET204_XI39/MM3717_g N_VSS_XI39/MM3717_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3625 XI39/NET4722 N_NET205_XI39/MM3625_g N_VSS_XI39/MM3625_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3640 N_NET482_XI39/MM3640_d N_NET206_XI39/MM3640_g N_VSS_XI39/MM3640_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3610 XI39/NET4782 N_NET207_XI39/MM3610_g N_VSS_XI39/MM3610_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3589 N_NET482_XI39/MM3589_d N_NET338_XI39/MM3589_g N_VSS_XI39/MM3589_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3674 XI39/NET6826 N_NET339_XI39/MM3674_g N_VSS_XI39/MM3674_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3653 N_NET482_XI39/MM3653_d N_NET340_XI39/MM3653_g N_VSS_XI39/MM3653_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3706 XI39/NET6698 N_NET211_XI39/MM3706_g N_VSS_XI39/MM3706_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3697 N_NET482_XI39/MM3697_d N_NET212_XI39/MM3697_g N_VSS_XI39/MM3697_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2730 XI39/NET8942 N_NET214_XI39/MM2730_g N_VSS_XI39/MM2730_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2745 N_NET482_XI39/MM2745_d N_NET215_XI39/MM2745_g N_VSS_XI39/MM2745_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2715 XI39/NET9002 N_NET216_XI39/MM2715_g N_VSS_XI39/MM2715_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2694 N_NET482_XI39/MM2694_d N_NET346_XI39/MM2694_g N_VSS_XI39/MM2694_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2779 XI39/NET8750 N_NET347_XI39/MM2779_g N_VSS_XI39/MM2779_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2758 N_NET482_XI39/MM2758_d N_NET348_XI39/MM2758_g N_VSS_XI39/MM2758_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2794 XI39/NET8690 N_NET349_XI39/MM2794_g N_VSS_XI39/MM2794_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2809 N_NET482_XI39/MM2809_d N_NET350_XI39/MM2809_g N_VSS_XI39/MM2809_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2651 XI39/NET9258 N_NET351_XI39/MM2651_g N_VSS_XI39/MM2651_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2630 N_NET482_XI39/MM2630_d N_NET352_XI39/MM2630_g N_VSS_XI39/MM2630_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2666 XI39/NET9198 N_NET224_XI39/MM2666_g N_VSS_XI39/MM2666_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2681 N_NET482_XI39/MM2681_d N_NET225_XI39/MM2681_g N_VSS_XI39/MM2681_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2602 XI39/NET9454 N_NET226_XI39/MM2602_g N_VSS_XI39/MM2602_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2617 N_NET482_XI39/MM2617_d N_NET356_XI39/MM2617_g N_VSS_XI39/MM2617_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2587 XI39/NET9514 N_NET357_XI39/MM2587_g N_VSS_XI39/MM2587_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2566 N_NET482_XI39/MM2566_d N_NET358_XI39/MM2566_g N_VSS_XI39/MM2566_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2907 XI39/NET8238 N_NET230_XI39/MM2907_g N_VSS_XI39/MM2907_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2886 N_NET482_XI39/MM2886_d N_NET360_XI39/MM2886_g N_VSS_XI39/MM2886_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2922 XI39/NET8178 N_NET361_XI39/MM2922_g N_VSS_XI39/MM2922_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2937 N_NET482_XI39/MM2937_d N_NET233_XI39/MM2937_g N_VSS_XI39/MM2937_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2858 XI39/NET8434 N_NET234_XI39/MM2858_g N_VSS_XI39/MM2858_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2873 N_NET482_XI39/MM2873_d N_NET235_XI39/MM2873_g N_VSS_XI39/MM2873_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2843 XI39/NET8494 N_NET365_XI39/MM2843_g N_VSS_XI39/MM2843_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2822 N_NET482_XI39/MM2822_d N_NET366_XI39/MM2822_g N_VSS_XI39/MM2822_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2986 XI39/NET7922 N_NET367_XI39/MM2986_g N_VSS_XI39/MM2986_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3001 N_NET482_XI39/MM3001_d N_NET368_XI39/MM3001_g N_VSS_XI39/MM3001_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2971 XI39/NET7982 N_NET369_XI39/MM2971_g N_VSS_XI39/MM2971_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2950 N_NET482_XI39/MM2950_d N_NET370_XI39/MM2950_g N_VSS_XI39/MM2950_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3035 XI39/NET7726 N_NET371_XI39/MM3035_g N_VSS_XI39/MM3035_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3014 N_NET482_XI39/MM3014_d N_NET242_XI39/MM3014_g N_VSS_XI39/MM3014_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3050 XI39/NET7666 N_NET373_XI39/MM3050_g N_VSS_XI39/MM3050_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3065 N_NET482_XI39/MM3065_d N_NET244_XI39/MM3065_g N_VSS_XI39/MM3065_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2389 XI39/NET10666 N_NET375_XI39/MM2389_g N_VSS_XI39/MM2389_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2374 N_NET482_XI39/MM2374_d N_NET376_XI39/MM2374_g N_VSS_XI39/MM2374_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2410 XI39/NET11230 N_NET377_XI39/MM2410_g N_VSS_XI39/MM2410_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2425 N_NET482_XI39/MM2425_d N_NET378_XI39/MM2425_g N_VSS_XI39/MM2425_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2346 XI39/NET10838 N_NET379_XI39/MM2346_g N_VSS_XI39/MM2346_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2361 N_NET482_XI39/MM2361_d N_NET380_XI39/MM2361_g N_VSS_XI39/MM2361_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2331 XI39/NET10898 N_NET381_XI39/MM2331_g N_VSS_XI39/MM2331_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2310 N_NET482_XI39/MM2310_d N_NET382_XI39/MM2310_g N_VSS_XI39/MM2310_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2476 XI39/NET11542 N_NET383_XI39/MM2476_g N_VSS_XI39/MM2476_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2489 N_NET482_XI39/MM2489_d N_NET384_XI39/MM2489_g N_VSS_XI39/MM2489_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2459 XI39/NET11034 N_NET385_XI39/MM2459_g N_VSS_XI39/MM2459_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2438 N_NET482_XI39/MM2438_d N_NET256_XI39/MM2438_g N_VSS_XI39/MM2438_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2523 XI39/NET11354 N_NET387_XI39/MM2523_g N_VSS_XI39/MM2523_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2502 N_NET482_XI39/MM2502_d N_NET388_XI39/MM2502_g N_VSS_XI39/MM2502_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2532 XI39/NET11318 N_NET389_XI39/MM2532_g N_VSS_XI39/MM2532_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2553 N_NET482_XI39/MM2553_d N_NET390_XI39/MM2553_g N_VSS_XI39/MM2553_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2218 XI39/NET10478 N_NET391_XI39/MM2218_g N_VSS_XI39/MM2218_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2233 N_NET482_XI39/MM2233_d N_NET262_XI39/MM2233_g N_VSS_XI39/MM2233_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2203 XI39/NET10538 N_NET263_XI39/MM2203_g N_VSS_XI39/MM2203_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2182 N_NET482_XI39/MM2182_d N_NET264_XI39/MM2182_g N_VSS_XI39/MM2182_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2267 XI39/NET10290 N_NET265_XI39/MM2267_g N_VSS_XI39/MM2267_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2246 N_NET482_XI39/MM2246_d N_NET396_XI39/MM2246_g N_VSS_XI39/MM2246_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2282 XI39/NET10230 N_NET267_XI39/MM2282_g N_VSS_XI39/MM2282_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2297 N_NET482_XI39/MM2297_d N_NET268_XI39/MM2297_g N_VSS_XI39/MM2297_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2133 XI39/NET9798 N_NET269_XI39/MM2133_g N_VSS_XI39/MM2133_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2118 N_NET482_XI39/MM2118_d N_NET270_XI39/MM2118_g N_VSS_XI39/MM2118_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2154 XI39/NET9714 N_NET401_XI39/MM2154_g N_VSS_XI39/MM2154_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2169 N_NET482_XI39/MM2169_d N_NET272_XI39/MM2169_g N_VSS_XI39/MM2169_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2090 XI39/NET9966 N_NET273_XI39/MM2090_g N_VSS_XI39/MM2090_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2105 N_NET482_XI39/MM2105_d N_NET404_XI39/MM2105_g N_VSS_XI39/MM2105_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2069 XI39/NET10026 N_NET405_XI39/MM2069_g N_VSS_XI39/MM2069_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM9 N_NET482_XI39/MM9_d N_NET0390_XI39/MM9_g N_VSS_XI39/MM9_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI54/XI1/XI8/XI3/MM2 N_XI54/XI1/XI8/NET12_XI54/XI1/XI8/XI3/MM2_d
+ N_NET068_XI54/XI1/XI8/XI3/MM2_g
+ N_XI54/XI1/XI8/XI3/NET13_XI54/XI1/XI8/XI3/MM2_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.3265e-13
+ AS=1.68025e-13 PD=1.46e-06 PS=7.15e-07
mXI54/XI1/XI7/XI3/MM2 N_XI54/XI1/XI7/NET12_XI54/XI1/XI7/XI3/MM2_d
+ N_NET068_XI54/XI1/XI7/XI3/MM2_g
+ N_XI54/XI1/XI7/XI3/NET13_XI54/XI1/XI7/XI3/MM2_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.3265e-13
+ AS=1.68025e-13 PD=1.46e-06 PS=7.15e-07
mXI29/XI1/MM41 N_NET420_XI29/XI1/MM41_d N_XI29/XI1/NET223_XI29/XI1/MM41_g
+ N_NET065_XI29/XI1/MM41_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI29/XI1/XI10/MM1 N_XI29/XI1/NET223_XI29/XI1/XI10/MM1_d
+ N_NET468_XI29/XI1/XI10/MM1_g N_VSS_XI29/XI1/XI10/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI29/XI1/MM42 N_NET421_XI29/XI1/MM42_d N_XI29/XI1/NET215_XI29/XI1/MM42_g
+ N_NET065_XI29/XI1/MM42_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI29/XI1/XI11/MM1 N_XI29/XI1/NET215_XI29/XI1/XI11/MM1_d
+ N_NET467_XI29/XI1/XI11/MM1_g N_VSS_XI29/XI1/XI11/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI39/MM3417 N_NET420_XI39/MM3417_d N_NET0133_XI39/MM3417_g N_VSS_XI39/MM3417_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3401 XI39/NET5618 N_NET280_XI39/MM3401_g N_VSS_XI39/MM3401_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3428 N_NET420_XI39/MM3428_d N_NET281_XI39/MM3428_g N_VSS_XI39/MM3428_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3447 XI39/NET5434 N_NET282_XI39/MM3447_g N_VSS_XI39/MM3447_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3365 N_NET420_XI39/MM3365_d N_NET153_XI39/MM3365_g N_VSS_XI39/MM3365_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3384 XI39/NET5686 N_NET284_XI39/MM3384_g N_VSS_XI39/MM3384_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3354 N_NET420_XI39/MM3354_d N_NET285_XI39/MM3354_g N_VSS_XI39/MM3354_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3333 XI39/NET3590 N_NET286_XI39/MM3333_g N_VSS_XI39/MM3333_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3492 N_NET420_XI39/MM3492_d N_NET287_XI39/MM3492_g N_VSS_XI39/MM3492_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3511 XI39/NET5178 N_NET158_XI39/MM3511_g N_VSS_XI39/MM3511_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3481 N_NET420_XI39/MM3481_d N_NET159_XI39/MM3481_g N_VSS_XI39/MM3481_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3464 XI39/NET5366 N_NET160_XI39/MM3464_g N_VSS_XI39/MM3464_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3545 N_NET420_XI39/MM3545_d N_NET291_XI39/MM3545_g N_VSS_XI39/MM3545_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3528 XI39/NET5110 N_NET162_XI39/MM3528_g N_VSS_XI39/MM3528_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3556 N_NET420_XI39/MM3556_d N_NET293_XI39/MM3556_g N_VSS_XI39/MM3556_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3575 XI39/NET4922 N_NET294_XI39/MM3575_g N_VSS_XI39/MM3575_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3237 N_NET420_XI39/MM3237_d N_NET295_XI39/MM3237_g N_VSS_XI39/MM3237_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3256 XI39/NET3898 N_NET296_XI39/MM3256_g N_VSS_XI39/MM3256_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3226 N_NET420_XI39/MM3226_d N_NET297_XI39/MM3226_g N_VSS_XI39/MM3226_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3209 XI39/NET4086 N_NET298_XI39/MM3209_g N_VSS_XI39/MM3209_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3290 N_NET420_XI39/MM3290_d N_NET299_XI39/MM3290_g N_VSS_XI39/MM3290_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3273 XI39/NET3830 N_NET170_XI39/MM3273_g N_VSS_XI39/MM3273_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3301 N_NET420_XI39/MM3301_d N_NET171_XI39/MM3301_g N_VSS_XI39/MM3301_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3320 XI39/NET3642 N_NET172_XI39/MM3320_g N_VSS_XI39/MM3320_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3162 N_NET420_XI39/MM3162_d N_NET303_XI39/MM3162_g N_VSS_XI39/MM3162_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3145 XI39/NET4342 N_NET304_XI39/MM3145_g N_VSS_XI39/MM3145_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3173 N_NET420_XI39/MM3173_d N_NET305_XI39/MM3173_g N_VSS_XI39/MM3173_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3192 XI39/NET4154 N_NET306_XI39/MM3192_g N_VSS_XI39/MM3192_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3109 N_NET420_XI39/MM3109_d N_NET307_XI39/MM3109_g N_VSS_XI39/MM3109_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3128 XI39/NET4410 N_NET308_XI39/MM3128_g N_VSS_XI39/MM3128_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3098 N_NET420_XI39/MM3098_d N_NET309_XI39/MM3098_g N_VSS_XI39/MM3098_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3081 XI39/NET4598 N_NET310_XI39/MM3081_g N_VSS_XI39/MM3081_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4000 N_NET420_XI39/MM4000_d N_NET311_XI39/MM4000_g N_VSS_XI39/MM4000_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3857 XI39/NET6094 N_NET312_XI39/MM3857_g N_VSS_XI39/MM3857_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3989 N_NET420_XI39/MM3989_d N_NET313_XI39/MM3989_g N_VSS_XI39/MM3989_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3972 XI39/NET7430 N_NET314_XI39/MM3972_g N_VSS_XI39/MM3972_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3891 N_NET420_XI39/MM3891_d N_NET315_XI39/MM3891_g N_VSS_XI39/MM3891_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3874 XI39/NET6026 N_NET316_XI39/MM3874_g N_VSS_XI39/MM3874_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3902 N_NET420_XI39/MM3902_d N_NET317_XI39/MM3902_g N_VSS_XI39/MM3902_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3921 XI39/NET5838 N_NET318_XI39/MM3921_g N_VSS_XI39/MM3921_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4069 N_NET420_XI39/MM4069_d N_NET319_XI39/MM4069_g N_VSS_XI39/MM4069_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4052 XI39/NET7110 N_NET320_XI39/MM4052_g N_VSS_XI39/MM4052_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3936 N_NET420_XI39/MM3936_d N_NET321_XI39/MM3936_g N_VSS_XI39/MM3936_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3955 XI39/NET7498 N_NET192_XI39/MM3955_g N_VSS_XI39/MM3955_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4016 N_NET420_XI39/MM4016_d N_NET193_XI39/MM4016_g N_VSS_XI39/MM4016_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4035 XI39/NET7178 N_NET194_XI39/MM4035_g N_VSS_XI39/MM4035_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4005 N_NET420_XI39/MM4005_d N_NET195_XI39/MM4005_g N_VSS_XI39/MM4005_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4082 XI39/NET6990 N_NET196_XI39/MM4082_g N_VSS_XI39/MM4082_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3801 N_NET420_XI39/MM3801_d N_NET197_XI39/MM3801_g N_VSS_XI39/MM3801_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3784 XI39/NET6386 N_NET198_XI39/MM3784_g N_VSS_XI39/MM3784_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3812 N_NET420_XI39/MM3812_d N_NET199_XI39/MM3812_g N_VSS_XI39/MM3812_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3831 XI39/NET6198 N_NET200_XI39/MM3831_g N_VSS_XI39/MM3831_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3748 N_NET420_XI39/MM3748_d N_NET331_XI39/MM3748_g N_VSS_XI39/MM3748_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3767 XI39/NET6454 N_NET332_XI39/MM3767_g N_VSS_XI39/MM3767_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3737 N_NET420_XI39/MM3737_d N_NET203_XI39/MM3737_g N_VSS_XI39/MM3737_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3720 XI39/NET6642 N_NET204_XI39/MM3720_g N_VSS_XI39/MM3720_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3620 N_NET420_XI39/MM3620_d N_NET205_XI39/MM3620_g N_VSS_XI39/MM3620_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3639 XI39/NET4666 N_NET206_XI39/MM3639_g N_VSS_XI39/MM3639_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3609 N_NET420_XI39/MM3609_d N_NET207_XI39/MM3609_g N_VSS_XI39/MM3609_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3592 XI39/NET4854 N_NET338_XI39/MM3592_g N_VSS_XI39/MM3592_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3673 N_NET420_XI39/MM3673_d N_NET339_XI39/MM3673_g N_VSS_XI39/MM3673_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3656 XI39/NET6898 N_NET340_XI39/MM3656_g N_VSS_XI39/MM3656_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3705 N_NET420_XI39/MM3705_d N_NET211_XI39/MM3705_g N_VSS_XI39/MM3705_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3696 XI39/NET6738 N_NET212_XI39/MM3696_g N_VSS_XI39/MM3696_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2725 N_NET420_XI39/MM2725_d N_NET214_XI39/MM2725_g N_VSS_XI39/MM2725_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2744 XI39/NET8890 N_NET215_XI39/MM2744_g N_VSS_XI39/MM2744_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2714 N_NET420_XI39/MM2714_d N_NET216_XI39/MM2714_g N_VSS_XI39/MM2714_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2697 XI39/NET9074 N_NET346_XI39/MM2697_g N_VSS_XI39/MM2697_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2778 N_NET420_XI39/MM2778_d N_NET347_XI39/MM2778_g N_VSS_XI39/MM2778_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2761 XI39/NET8822 N_NET348_XI39/MM2761_g N_VSS_XI39/MM2761_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2789 N_NET420_XI39/MM2789_d N_NET349_XI39/MM2789_g N_VSS_XI39/MM2789_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2808 XI39/NET8634 N_NET350_XI39/MM2808_g N_VSS_XI39/MM2808_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2650 N_NET420_XI39/MM2650_d N_NET351_XI39/MM2650_g N_VSS_XI39/MM2650_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2633 XI39/NET9330 N_NET352_XI39/MM2633_g N_VSS_XI39/MM2633_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2661 N_NET420_XI39/MM2661_d N_NET224_XI39/MM2661_g N_VSS_XI39/MM2661_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2680 XI39/NET9142 N_NET225_XI39/MM2680_g N_VSS_XI39/MM2680_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2597 N_NET420_XI39/MM2597_d N_NET226_XI39/MM2597_g N_VSS_XI39/MM2597_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2616 XI39/NET9398 N_NET356_XI39/MM2616_g N_VSS_XI39/MM2616_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2586 N_NET420_XI39/MM2586_d N_NET357_XI39/MM2586_g N_VSS_XI39/MM2586_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2569 XI39/NET9586 N_NET358_XI39/MM2569_g N_VSS_XI39/MM2569_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2906 N_NET420_XI39/MM2906_d N_NET230_XI39/MM2906_g N_VSS_XI39/MM2906_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2889 XI39/NET8310 N_NET360_XI39/MM2889_g N_VSS_XI39/MM2889_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2917 N_NET420_XI39/MM2917_d N_NET361_XI39/MM2917_g N_VSS_XI39/MM2917_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2936 XI39/NET8122 N_NET233_XI39/MM2936_g N_VSS_XI39/MM2936_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2853 N_NET420_XI39/MM2853_d N_NET234_XI39/MM2853_g N_VSS_XI39/MM2853_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2872 XI39/NET8378 N_NET235_XI39/MM2872_g N_VSS_XI39/MM2872_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2842 N_NET420_XI39/MM2842_d N_NET365_XI39/MM2842_g N_VSS_XI39/MM2842_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2825 XI39/NET8566 N_NET366_XI39/MM2825_g N_VSS_XI39/MM2825_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2981 N_NET420_XI39/MM2981_d N_NET367_XI39/MM2981_g N_VSS_XI39/MM2981_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3000 XI39/NET7866 N_NET368_XI39/MM3000_g N_VSS_XI39/MM3000_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2970 N_NET420_XI39/MM2970_d N_NET369_XI39/MM2970_g N_VSS_XI39/MM2970_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2953 XI39/NET8054 N_NET370_XI39/MM2953_g N_VSS_XI39/MM2953_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3034 N_NET420_XI39/MM3034_d N_NET371_XI39/MM3034_g N_VSS_XI39/MM3034_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3017 XI39/NET7798 N_NET242_XI39/MM3017_g N_VSS_XI39/MM3017_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3045 N_NET420_XI39/MM3045_d N_NET373_XI39/MM3045_g N_VSS_XI39/MM3045_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3064 XI39/NET7610 N_NET244_XI39/MM3064_g N_VSS_XI39/MM3064_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2394 N_NET420_XI39/MM2394_d N_NET375_XI39/MM2394_g N_VSS_XI39/MM2394_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2377 XI39/NET10714 N_NET376_XI39/MM2377_g N_VSS_XI39/MM2377_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2405 N_NET420_XI39/MM2405_d N_NET377_XI39/MM2405_g N_VSS_XI39/MM2405_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2424 XI39/NET11174 N_NET378_XI39/MM2424_g N_VSS_XI39/MM2424_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2341 N_NET420_XI39/MM2341_d N_NET379_XI39/MM2341_g N_VSS_XI39/MM2341_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2360 XI39/NET10782 N_NET380_XI39/MM2360_g N_VSS_XI39/MM2360_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2330 N_NET420_XI39/MM2330_d N_NET381_XI39/MM2330_g N_VSS_XI39/MM2330_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2313 XI39/NET10970 N_NET382_XI39/MM2313_g N_VSS_XI39/MM2313_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2469 N_NET420_XI39/MM2469_d N_NET383_XI39/MM2469_g N_VSS_XI39/MM2469_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2488 XI39/NET11494 N_NET384_XI39/MM2488_g N_VSS_XI39/MM2488_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2458 N_NET420_XI39/MM2458_d N_NET385_XI39/MM2458_g N_VSS_XI39/MM2458_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2441 XI39/NET11106 N_NET256_XI39/MM2441_g N_VSS_XI39/MM2441_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2522 N_NET420_XI39/MM2522_d N_NET387_XI39/MM2522_g N_VSS_XI39/MM2522_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2505 XI39/NET11426 N_NET388_XI39/MM2505_g N_VSS_XI39/MM2505_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2533 N_NET420_XI39/MM2533_d N_NET389_XI39/MM2533_g N_VSS_XI39/MM2533_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2552 XI39/NET11614 N_NET390_XI39/MM2552_g N_VSS_XI39/MM2552_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2213 N_NET420_XI39/MM2213_d N_NET391_XI39/MM2213_g N_VSS_XI39/MM2213_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2232 XI39/NET10426 N_NET262_XI39/MM2232_g N_VSS_XI39/MM2232_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2202 N_NET420_XI39/MM2202_d N_NET263_XI39/MM2202_g N_VSS_XI39/MM2202_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2185 XI39/NET10606 N_NET264_XI39/MM2185_g N_VSS_XI39/MM2185_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2266 N_NET420_XI39/MM2266_d N_NET265_XI39/MM2266_g N_VSS_XI39/MM2266_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2249 XI39/NET10358 N_NET396_XI39/MM2249_g N_VSS_XI39/MM2249_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2277 N_NET420_XI39/MM2277_d N_NET267_XI39/MM2277_g N_VSS_XI39/MM2277_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2296 XI39/NET10178 N_NET268_XI39/MM2296_g N_VSS_XI39/MM2296_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2138 N_NET420_XI39/MM2138_d N_NET269_XI39/MM2138_g N_VSS_XI39/MM2138_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2121 XI39/NET9842 N_NET270_XI39/MM2121_g N_VSS_XI39/MM2121_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2149 N_NET420_XI39/MM2149_d N_NET401_XI39/MM2149_g N_VSS_XI39/MM2149_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2168 XI39/NET9662 N_NET272_XI39/MM2168_g N_VSS_XI39/MM2168_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2085 N_NET420_XI39/MM2085_d N_NET273_XI39/MM2085_g N_VSS_XI39/MM2085_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2104 XI39/NET9914 N_NET404_XI39/MM2104_g N_VSS_XI39/MM2104_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2074 N_NET420_XI39/MM2074_d N_NET405_XI39/MM2074_g N_VSS_XI39/MM2074_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2 XI39/NET10050 N_NET0390_XI39/MM2_g N_VSS_XI39/MM2_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3420 XI39/NET5542 N_NET0133_XI39/MM3420_g N_VSS_XI39/MM3420_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3396 N_NET421_XI39/MM3396_d N_NET280_XI39/MM3396_g N_VSS_XI39/MM3396_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3427 XI39/NET5514 N_NET281_XI39/MM3427_g N_VSS_XI39/MM3427_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3450 N_NET421_XI39/MM3450_d N_NET282_XI39/MM3450_g N_VSS_XI39/MM3450_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3364 XI39/NET5766 N_NET153_XI39/MM3364_g N_VSS_XI39/MM3364_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3387 N_NET421_XI39/MM3387_d N_NET284_XI39/MM3387_g N_VSS_XI39/MM3387_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3349 XI39/NET3526 N_NET285_XI39/MM3349_g N_VSS_XI39/MM3349_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3332 N_NET421_XI39/MM3332_d N_NET286_XI39/MM3332_g N_VSS_XI39/MM3332_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3491 XI39/NET5258 N_NET287_XI39/MM3491_g N_VSS_XI39/MM3491_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3514 N_NET421_XI39/MM3514_d N_NET158_XI39/MM3514_g N_VSS_XI39/MM3514_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3476 XI39/NET5318 N_NET159_XI39/MM3476_g N_VSS_XI39/MM3476_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3459 N_NET421_XI39/MM3459_d N_NET160_XI39/MM3459_g N_VSS_XI39/MM3459_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3540 XI39/NET5062 N_NET291_XI39/MM3540_g N_VSS_XI39/MM3540_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3523 N_NET421_XI39/MM3523_d N_NET162_XI39/MM3523_g N_VSS_XI39/MM3523_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3555 XI39/NET5002 N_NET293_XI39/MM3555_g N_VSS_XI39/MM3555_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3578 N_NET421_XI39/MM3578_d N_NET294_XI39/MM3578_g N_VSS_XI39/MM3578_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3236 XI39/NET3978 N_NET295_XI39/MM3236_g N_VSS_XI39/MM3236_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3259 N_NET421_XI39/MM3259_d N_NET296_XI39/MM3259_g N_VSS_XI39/MM3259_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3221 XI39/NET4038 N_NET297_XI39/MM3221_g N_VSS_XI39/MM3221_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3204 N_NET421_XI39/MM3204_d N_NET298_XI39/MM3204_g N_VSS_XI39/MM3204_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3285 XI39/NET3782 N_NET299_XI39/MM3285_g N_VSS_XI39/MM3285_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3268 N_NET421_XI39/MM3268_d N_NET170_XI39/MM3268_g N_VSS_XI39/MM3268_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3300 XI39/NET3722 N_NET171_XI39/MM3300_g N_VSS_XI39/MM3300_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3323 N_NET421_XI39/MM3323_d N_NET172_XI39/MM3323_g N_VSS_XI39/MM3323_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3157 XI39/NET4294 N_NET303_XI39/MM3157_g N_VSS_XI39/MM3157_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3140 N_NET421_XI39/MM3140_d N_NET304_XI39/MM3140_g N_VSS_XI39/MM3140_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3172 XI39/NET4234 N_NET305_XI39/MM3172_g N_VSS_XI39/MM3172_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3195 N_NET421_XI39/MM3195_d N_NET306_XI39/MM3195_g N_VSS_XI39/MM3195_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3108 XI39/NET4490 N_NET307_XI39/MM3108_g N_VSS_XI39/MM3108_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3131 N_NET421_XI39/MM3131_d N_NET308_XI39/MM3131_g N_VSS_XI39/MM3131_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3093 XI39/NET4550 N_NET309_XI39/MM3093_g N_VSS_XI39/MM3093_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3076 N_NET421_XI39/MM3076_d N_NET310_XI39/MM3076_g N_VSS_XI39/MM3076_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3999 XI39/NET7322 N_NET311_XI39/MM3999_g N_VSS_XI39/MM3999_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3860 N_NET421_XI39/MM3860_d N_NET312_XI39/MM3860_g N_VSS_XI39/MM3860_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3984 XI39/NET7382 N_NET313_XI39/MM3984_g N_VSS_XI39/MM3984_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3967 N_NET421_XI39/MM3967_d N_NET314_XI39/MM3967_g N_VSS_XI39/MM3967_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3886 XI39/NET5978 N_NET315_XI39/MM3886_g N_VSS_XI39/MM3886_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3869 N_NET421_XI39/MM3869_d N_NET316_XI39/MM3869_g N_VSS_XI39/MM3869_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3901 XI39/NET5918 N_NET317_XI39/MM3901_g N_VSS_XI39/MM3901_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3924 N_NET421_XI39/MM3924_d N_NET318_XI39/MM3924_g N_VSS_XI39/MM3924_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4064 XI39/NET7062 N_NET319_XI39/MM4064_g N_VSS_XI39/MM4064_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4047 N_NET421_XI39/MM4047_d N_NET320_XI39/MM4047_g N_VSS_XI39/MM4047_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3939 XI39/NET7562 N_NET321_XI39/MM3939_g N_VSS_XI39/MM3939_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3958 N_NET421_XI39/MM3958_d N_NET192_XI39/MM3958_g N_VSS_XI39/MM3958_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4015 XI39/NET7258 N_NET193_XI39/MM4015_g N_VSS_XI39/MM4015_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4038 N_NET421_XI39/MM4038_d N_NET194_XI39/MM4038_g N_VSS_XI39/MM4038_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4006 XI39/NET7294 N_NET195_XI39/MM4006_g N_VSS_XI39/MM4006_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4077 N_NET421_XI39/MM4077_d N_NET196_XI39/MM4077_g N_VSS_XI39/MM4077_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3796 XI39/NET6338 N_NET197_XI39/MM3796_g N_VSS_XI39/MM3796_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3779 N_NET421_XI39/MM3779_d N_NET198_XI39/MM3779_g N_VSS_XI39/MM3779_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3811 XI39/NET6278 N_NET199_XI39/MM3811_g N_VSS_XI39/MM3811_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3834 N_NET421_XI39/MM3834_d N_NET200_XI39/MM3834_g N_VSS_XI39/MM3834_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3747 XI39/NET6534 N_NET331_XI39/MM3747_g N_VSS_XI39/MM3747_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3770 N_NET421_XI39/MM3770_d N_NET332_XI39/MM3770_g N_VSS_XI39/MM3770_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3732 XI39/NET6594 N_NET203_XI39/MM3732_g N_VSS_XI39/MM3732_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3715 N_NET421_XI39/MM3715_d N_NET204_XI39/MM3715_g N_VSS_XI39/MM3715_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3619 XI39/NET4746 N_NET205_XI39/MM3619_g N_VSS_XI39/MM3619_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3642 N_NET421_XI39/MM3642_d N_NET206_XI39/MM3642_g N_VSS_XI39/MM3642_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3604 XI39/NET4806 N_NET207_XI39/MM3604_g N_VSS_XI39/MM3604_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3587 N_NET421_XI39/MM3587_d N_NET338_XI39/MM3587_g N_VSS_XI39/MM3587_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3668 XI39/NET6850 N_NET339_XI39/MM3668_g N_VSS_XI39/MM3668_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3651 N_NET421_XI39/MM3651_d N_NET340_XI39/MM3651_g N_VSS_XI39/MM3651_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3684 XI39/NET6786 N_NET211_XI39/MM3684_g N_VSS_XI39/MM3684_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3699 N_NET421_XI39/MM3699_d N_NET212_XI39/MM3699_g N_VSS_XI39/MM3699_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2724 XI39/NET8966 N_NET214_XI39/MM2724_g N_VSS_XI39/MM2724_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2747 N_NET421_XI39/MM2747_d N_NET215_XI39/MM2747_g N_VSS_XI39/MM2747_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2709 XI39/NET9026 N_NET216_XI39/MM2709_g N_VSS_XI39/MM2709_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2692 N_NET421_XI39/MM2692_d N_NET346_XI39/MM2692_g N_VSS_XI39/MM2692_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2773 XI39/NET8774 N_NET347_XI39/MM2773_g N_VSS_XI39/MM2773_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2756 N_NET421_XI39/MM2756_d N_NET348_XI39/MM2756_g N_VSS_XI39/MM2756_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2788 XI39/NET8714 N_NET349_XI39/MM2788_g N_VSS_XI39/MM2788_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2811 N_NET421_XI39/MM2811_d N_NET350_XI39/MM2811_g N_VSS_XI39/MM2811_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2645 XI39/NET9282 N_NET351_XI39/MM2645_g N_VSS_XI39/MM2645_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2628 N_NET421_XI39/MM2628_d N_NET352_XI39/MM2628_g N_VSS_XI39/MM2628_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2660 XI39/NET9222 N_NET224_XI39/MM2660_g N_VSS_XI39/MM2660_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2683 N_NET421_XI39/MM2683_d N_NET225_XI39/MM2683_g N_VSS_XI39/MM2683_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2596 XI39/NET9478 N_NET226_XI39/MM2596_g N_VSS_XI39/MM2596_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2619 N_NET421_XI39/MM2619_d N_NET356_XI39/MM2619_g N_VSS_XI39/MM2619_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2581 XI39/NET9538 N_NET357_XI39/MM2581_g N_VSS_XI39/MM2581_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2564 N_NET421_XI39/MM2564_d N_NET358_XI39/MM2564_g N_VSS_XI39/MM2564_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2901 XI39/NET8262 N_NET230_XI39/MM2901_g N_VSS_XI39/MM2901_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2884 N_NET421_XI39/MM2884_d N_NET360_XI39/MM2884_g N_VSS_XI39/MM2884_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2916 XI39/NET8202 N_NET361_XI39/MM2916_g N_VSS_XI39/MM2916_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2939 N_NET421_XI39/MM2939_d N_NET233_XI39/MM2939_g N_VSS_XI39/MM2939_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2852 XI39/NET8458 N_NET234_XI39/MM2852_g N_VSS_XI39/MM2852_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2875 N_NET421_XI39/MM2875_d N_NET235_XI39/MM2875_g N_VSS_XI39/MM2875_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2837 XI39/NET8518 N_NET365_XI39/MM2837_g N_VSS_XI39/MM2837_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2820 N_NET421_XI39/MM2820_d N_NET366_XI39/MM2820_g N_VSS_XI39/MM2820_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2980 XI39/NET7946 N_NET367_XI39/MM2980_g N_VSS_XI39/MM2980_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3003 N_NET421_XI39/MM3003_d N_NET368_XI39/MM3003_g N_VSS_XI39/MM3003_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2965 XI39/NET8006 N_NET369_XI39/MM2965_g N_VSS_XI39/MM2965_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2948 N_NET421_XI39/MM2948_d N_NET370_XI39/MM2948_g N_VSS_XI39/MM2948_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3029 XI39/NET7750 N_NET371_XI39/MM3029_g N_VSS_XI39/MM3029_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3012 N_NET421_XI39/MM3012_d N_NET242_XI39/MM3012_g N_VSS_XI39/MM3012_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3044 XI39/NET7690 N_NET373_XI39/MM3044_g N_VSS_XI39/MM3044_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3067 N_NET421_XI39/MM3067_d N_NET244_XI39/MM3067_g N_VSS_XI39/MM3067_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2399 XI39/NET11274 N_NET375_XI39/MM2399_g N_VSS_XI39/MM2399_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2372 N_NET421_XI39/MM2372_d N_NET376_XI39/MM2372_g N_VSS_XI39/MM2372_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2404 XI39/NET11254 N_NET377_XI39/MM2404_g N_VSS_XI39/MM2404_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2427 N_NET421_XI39/MM2427_d N_NET378_XI39/MM2427_g N_VSS_XI39/MM2427_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2340 XI39/NET10862 N_NET379_XI39/MM2340_g N_VSS_XI39/MM2340_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2363 N_NET421_XI39/MM2363_d N_NET380_XI39/MM2363_g N_VSS_XI39/MM2363_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2325 XI39/NET10922 N_NET381_XI39/MM2325_g N_VSS_XI39/MM2325_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2308 N_NET421_XI39/MM2308_d N_NET382_XI39/MM2308_g N_VSS_XI39/MM2308_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2470 XI39/NET11566 N_NET383_XI39/MM2470_g N_VSS_XI39/MM2470_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2491 N_NET421_XI39/MM2491_d N_NET384_XI39/MM2491_g N_VSS_XI39/MM2491_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2453 XI39/NET11058 N_NET385_XI39/MM2453_g N_VSS_XI39/MM2453_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2436 N_NET421_XI39/MM2436_d N_NET256_XI39/MM2436_g N_VSS_XI39/MM2436_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2517 XI39/NET11378 N_NET387_XI39/MM2517_g N_VSS_XI39/MM2517_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2500 N_NET421_XI39/MM2500_d N_NET388_XI39/MM2500_g N_VSS_XI39/MM2500_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2542 XI39/NET11654 N_NET389_XI39/MM2542_g N_VSS_XI39/MM2542_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2555 N_NET421_XI39/MM2555_d N_NET390_XI39/MM2555_g N_VSS_XI39/MM2555_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2212 XI39/NET10502 N_NET391_XI39/MM2212_g N_VSS_XI39/MM2212_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2235 N_NET421_XI39/MM2235_d N_NET262_XI39/MM2235_g N_VSS_XI39/MM2235_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2197 XI39/NET10562 N_NET263_XI39/MM2197_g N_VSS_XI39/MM2197_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2180 N_NET421_XI39/MM2180_d N_NET264_XI39/MM2180_g N_VSS_XI39/MM2180_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2261 XI39/NET10314 N_NET265_XI39/MM2261_g N_VSS_XI39/MM2261_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2244 N_NET421_XI39/MM2244_d N_NET396_XI39/MM2244_g N_VSS_XI39/MM2244_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2276 XI39/NET10254 N_NET267_XI39/MM2276_g N_VSS_XI39/MM2276_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2299 N_NET421_XI39/MM2299_d N_NET268_XI39/MM2299_g N_VSS_XI39/MM2299_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2141 XI39/NET9766 N_NET269_XI39/MM2141_g N_VSS_XI39/MM2141_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2116 N_NET421_XI39/MM2116_d N_NET270_XI39/MM2116_g N_VSS_XI39/MM2116_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2148 XI39/NET9738 N_NET401_XI39/MM2148_g N_VSS_XI39/MM2148_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2171 N_NET421_XI39/MM2171_d N_NET272_XI39/MM2171_g N_VSS_XI39/MM2171_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2084 XI39/NET9990 N_NET273_XI39/MM2084_g N_VSS_XI39/MM2084_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2107 N_NET421_XI39/MM2107_d N_NET404_XI39/MM2107_g N_VSS_XI39/MM2107_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2075 XI39/NET10114 N_NET405_XI39/MM2075_g N_VSS_XI39/MM2075_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM11 N_NET421_XI39/MM11_d N_NET0390_XI39/MM11_g N_VSS_XI39/MM11_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI54/XI1/XI8/XI2/MM1 N_XI54/XI1/NET9_XI54/XI1/XI8/XI2/MM1_d
+ N_XI54/XI1/XI8/NET12_XI54/XI1/XI8/XI2/MM1_g N_VSS_XI54/XI1/XI8/XI2/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13
+ AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI54/XI1/XI7/XI2/MM1 N_XI54/XI1/NET10_XI54/XI1/XI7/XI2/MM1_d
+ N_XI54/XI1/XI7/NET12_XI54/XI1/XI7/XI2/MM1_g N_VSS_XI54/XI1/XI7/XI2/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13
+ AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI29/XI1/MM43 N_NET485_XI29/XI1/MM43_d N_XI29/XI1/NET211_XI29/XI1/MM43_g
+ N_NET065_XI29/XI1/MM43_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI29/XI1/XI12/MM1 N_XI29/XI1/NET211_XI29/XI1/XI12/MM1_d
+ N_NET466_XI29/XI1/XI12/MM1_g N_VSS_XI29/XI1/XI12/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI29/XI1/MM44 N_NET486_XI29/XI1/MM44_d N_XI29/XI1/NET203_XI29/XI1/MM44_g
+ N_NET065_XI29/XI1/MM44_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI29/XI1/XI13/MM1 N_XI29/XI1/NET203_XI29/XI1/XI13/MM1_d
+ N_NET465_XI29/XI1/XI13/MM1_g N_VSS_XI29/XI1/XI13/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI39/MM3419 N_NET485_XI39/MM3419_d N_NET0133_XI39/MM3419_g N_VSS_XI39/MM3419_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3403 XI39/NET5610 N_NET280_XI39/MM3403_g N_VSS_XI39/MM3403_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3426 N_NET485_XI39/MM3426_d N_NET281_XI39/MM3426_g N_VSS_XI39/MM3426_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3449 XI39/NET5426 N_NET282_XI39/MM3449_g N_VSS_XI39/MM3449_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3363 N_NET485_XI39/MM3363_d N_NET153_XI39/MM3363_g N_VSS_XI39/MM3363_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3386 XI39/NET5678 N_NET284_XI39/MM3386_g N_VSS_XI39/MM3386_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3356 N_NET485_XI39/MM3356_d N_NET285_XI39/MM3356_g N_VSS_XI39/MM3356_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3331 XI39/NET3598 N_NET286_XI39/MM3331_g N_VSS_XI39/MM3331_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3490 N_NET485_XI39/MM3490_d N_NET287_XI39/MM3490_g N_VSS_XI39/MM3490_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3513 XI39/NET5170 N_NET158_XI39/MM3513_g N_VSS_XI39/MM3513_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3483 N_NET485_XI39/MM3483_d N_NET159_XI39/MM3483_g N_VSS_XI39/MM3483_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3466 XI39/NET5358 N_NET160_XI39/MM3466_g N_VSS_XI39/MM3466_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3547 N_NET485_XI39/MM3547_d N_NET291_XI39/MM3547_g N_VSS_XI39/MM3547_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3530 XI39/NET5102 N_NET162_XI39/MM3530_g N_VSS_XI39/MM3530_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3554 N_NET485_XI39/MM3554_d N_NET293_XI39/MM3554_g N_VSS_XI39/MM3554_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3577 XI39/NET4914 N_NET294_XI39/MM3577_g N_VSS_XI39/MM3577_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3235 N_NET485_XI39/MM3235_d N_NET295_XI39/MM3235_g N_VSS_XI39/MM3235_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3258 XI39/NET3890 N_NET296_XI39/MM3258_g N_VSS_XI39/MM3258_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3228 N_NET485_XI39/MM3228_d N_NET297_XI39/MM3228_g N_VSS_XI39/MM3228_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3211 XI39/NET4078 N_NET298_XI39/MM3211_g N_VSS_XI39/MM3211_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3292 N_NET485_XI39/MM3292_d N_NET299_XI39/MM3292_g N_VSS_XI39/MM3292_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3275 XI39/NET3822 N_NET170_XI39/MM3275_g N_VSS_XI39/MM3275_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3299 N_NET485_XI39/MM3299_d N_NET171_XI39/MM3299_g N_VSS_XI39/MM3299_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3322 XI39/NET3634 N_NET172_XI39/MM3322_g N_VSS_XI39/MM3322_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3164 N_NET485_XI39/MM3164_d N_NET303_XI39/MM3164_g N_VSS_XI39/MM3164_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3147 XI39/NET4334 N_NET304_XI39/MM3147_g N_VSS_XI39/MM3147_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3171 N_NET485_XI39/MM3171_d N_NET305_XI39/MM3171_g N_VSS_XI39/MM3171_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3194 XI39/NET4146 N_NET306_XI39/MM3194_g N_VSS_XI39/MM3194_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3107 N_NET485_XI39/MM3107_d N_NET307_XI39/MM3107_g N_VSS_XI39/MM3107_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3130 XI39/NET4402 N_NET308_XI39/MM3130_g N_VSS_XI39/MM3130_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3100 N_NET485_XI39/MM3100_d N_NET309_XI39/MM3100_g N_VSS_XI39/MM3100_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3083 XI39/NET4590 N_NET310_XI39/MM3083_g N_VSS_XI39/MM3083_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3998 N_NET485_XI39/MM3998_d N_NET311_XI39/MM3998_g N_VSS_XI39/MM3998_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3859 XI39/NET6086 N_NET312_XI39/MM3859_g N_VSS_XI39/MM3859_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3991 N_NET485_XI39/MM3991_d N_NET313_XI39/MM3991_g N_VSS_XI39/MM3991_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3974 XI39/NET7422 N_NET314_XI39/MM3974_g N_VSS_XI39/MM3974_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3893 N_NET485_XI39/MM3893_d N_NET315_XI39/MM3893_g N_VSS_XI39/MM3893_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3876 XI39/NET6018 N_NET316_XI39/MM3876_g N_VSS_XI39/MM3876_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3900 N_NET485_XI39/MM3900_d N_NET317_XI39/MM3900_g N_VSS_XI39/MM3900_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3923 XI39/NET5830 N_NET318_XI39/MM3923_g N_VSS_XI39/MM3923_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4071 N_NET485_XI39/MM4071_d N_NET319_XI39/MM4071_g N_VSS_XI39/MM4071_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4054 XI39/NET7102 N_NET320_XI39/MM4054_g N_VSS_XI39/MM4054_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3934 N_NET485_XI39/MM3934_d N_NET321_XI39/MM3934_g N_VSS_XI39/MM3934_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3957 XI39/NET7490 N_NET192_XI39/MM3957_g N_VSS_XI39/MM3957_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4014 N_NET485_XI39/MM4014_d N_NET193_XI39/MM4014_g N_VSS_XI39/MM4014_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4037 XI39/NET7170 N_NET194_XI39/MM4037_g N_VSS_XI39/MM4037_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4007 N_NET485_XI39/MM4007_d N_NET195_XI39/MM4007_g N_VSS_XI39/MM4007_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4084 XI39/NET6982 N_NET196_XI39/MM4084_g N_VSS_XI39/MM4084_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3803 N_NET485_XI39/MM3803_d N_NET197_XI39/MM3803_g N_VSS_XI39/MM3803_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3786 XI39/NET6378 N_NET198_XI39/MM3786_g N_VSS_XI39/MM3786_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3810 N_NET485_XI39/MM3810_d N_NET199_XI39/MM3810_g N_VSS_XI39/MM3810_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3833 XI39/NET6190 N_NET200_XI39/MM3833_g N_VSS_XI39/MM3833_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3746 N_NET485_XI39/MM3746_d N_NET331_XI39/MM3746_g N_VSS_XI39/MM3746_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3769 XI39/NET6446 N_NET332_XI39/MM3769_g N_VSS_XI39/MM3769_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3739 N_NET485_XI39/MM3739_d N_NET203_XI39/MM3739_g N_VSS_XI39/MM3739_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3722 XI39/NET6634 N_NET204_XI39/MM3722_g N_VSS_XI39/MM3722_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3618 N_NET485_XI39/MM3618_d N_NET205_XI39/MM3618_g N_VSS_XI39/MM3618_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3641 XI39/NET4658 N_NET206_XI39/MM3641_g N_VSS_XI39/MM3641_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3611 N_NET485_XI39/MM3611_d N_NET207_XI39/MM3611_g N_VSS_XI39/MM3611_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3594 XI39/NET4846 N_NET338_XI39/MM3594_g N_VSS_XI39/MM3594_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3675 N_NET485_XI39/MM3675_d N_NET339_XI39/MM3675_g N_VSS_XI39/MM3675_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3658 XI39/NET6890 N_NET340_XI39/MM3658_g N_VSS_XI39/MM3658_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3707 N_NET485_XI39/MM3707_d N_NET211_XI39/MM3707_g N_VSS_XI39/MM3707_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3698 XI39/NET6730 N_NET212_XI39/MM3698_g N_VSS_XI39/MM3698_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2723 N_NET485_XI39/MM2723_d N_NET214_XI39/MM2723_g N_VSS_XI39/MM2723_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2746 XI39/NET8882 N_NET215_XI39/MM2746_g N_VSS_XI39/MM2746_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2716 N_NET485_XI39/MM2716_d N_NET216_XI39/MM2716_g N_VSS_XI39/MM2716_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2699 XI39/NET9066 N_NET346_XI39/MM2699_g N_VSS_XI39/MM2699_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2780 N_NET485_XI39/MM2780_d N_NET347_XI39/MM2780_g N_VSS_XI39/MM2780_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2763 XI39/NET8814 N_NET348_XI39/MM2763_g N_VSS_XI39/MM2763_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2787 N_NET485_XI39/MM2787_d N_NET349_XI39/MM2787_g N_VSS_XI39/MM2787_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2810 XI39/NET8626 N_NET350_XI39/MM2810_g N_VSS_XI39/MM2810_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2652 N_NET485_XI39/MM2652_d N_NET351_XI39/MM2652_g N_VSS_XI39/MM2652_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2635 XI39/NET9322 N_NET352_XI39/MM2635_g N_VSS_XI39/MM2635_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2659 N_NET485_XI39/MM2659_d N_NET224_XI39/MM2659_g N_VSS_XI39/MM2659_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2682 XI39/NET9134 N_NET225_XI39/MM2682_g N_VSS_XI39/MM2682_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2595 N_NET485_XI39/MM2595_d N_NET226_XI39/MM2595_g N_VSS_XI39/MM2595_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2618 XI39/NET9390 N_NET356_XI39/MM2618_g N_VSS_XI39/MM2618_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2588 N_NET485_XI39/MM2588_d N_NET357_XI39/MM2588_g N_VSS_XI39/MM2588_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2571 XI39/NET9578 N_NET358_XI39/MM2571_g N_VSS_XI39/MM2571_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2908 N_NET485_XI39/MM2908_d N_NET230_XI39/MM2908_g N_VSS_XI39/MM2908_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2891 XI39/NET8302 N_NET360_XI39/MM2891_g N_VSS_XI39/MM2891_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2915 N_NET485_XI39/MM2915_d N_NET361_XI39/MM2915_g N_VSS_XI39/MM2915_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2938 XI39/NET8114 N_NET233_XI39/MM2938_g N_VSS_XI39/MM2938_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2851 N_NET485_XI39/MM2851_d N_NET234_XI39/MM2851_g N_VSS_XI39/MM2851_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2874 XI39/NET8370 N_NET235_XI39/MM2874_g N_VSS_XI39/MM2874_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2844 N_NET485_XI39/MM2844_d N_NET365_XI39/MM2844_g N_VSS_XI39/MM2844_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2827 XI39/NET8558 N_NET366_XI39/MM2827_g N_VSS_XI39/MM2827_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2979 N_NET485_XI39/MM2979_d N_NET367_XI39/MM2979_g N_VSS_XI39/MM2979_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3002 XI39/NET7858 N_NET368_XI39/MM3002_g N_VSS_XI39/MM3002_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2972 N_NET485_XI39/MM2972_d N_NET369_XI39/MM2972_g N_VSS_XI39/MM2972_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2955 XI39/NET8046 N_NET370_XI39/MM2955_g N_VSS_XI39/MM2955_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3036 N_NET485_XI39/MM3036_d N_NET371_XI39/MM3036_g N_VSS_XI39/MM3036_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3019 XI39/NET7790 N_NET242_XI39/MM3019_g N_VSS_XI39/MM3019_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3043 N_NET485_XI39/MM3043_d N_NET373_XI39/MM3043_g N_VSS_XI39/MM3043_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3066 XI39/NET7602 N_NET244_XI39/MM3066_g N_VSS_XI39/MM3066_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2396 N_NET485_XI39/MM2396_d N_NET375_XI39/MM2396_g N_VSS_XI39/MM2396_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2379 XI39/NET10706 N_NET376_XI39/MM2379_g N_VSS_XI39/MM2379_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2403 N_NET485_XI39/MM2403_d N_NET377_XI39/MM2403_g N_VSS_XI39/MM2403_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2426 XI39/NET11166 N_NET378_XI39/MM2426_g N_VSS_XI39/MM2426_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2339 N_NET485_XI39/MM2339_d N_NET379_XI39/MM2339_g N_VSS_XI39/MM2339_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2362 XI39/NET10774 N_NET380_XI39/MM2362_g N_VSS_XI39/MM2362_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2332 N_NET485_XI39/MM2332_d N_NET381_XI39/MM2332_g N_VSS_XI39/MM2332_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2315 XI39/NET10962 N_NET382_XI39/MM2315_g N_VSS_XI39/MM2315_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2467 N_NET485_XI39/MM2467_d N_NET383_XI39/MM2467_g N_VSS_XI39/MM2467_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2490 XI39/NET11486 N_NET384_XI39/MM2490_g N_VSS_XI39/MM2490_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2460 N_NET485_XI39/MM2460_d N_NET385_XI39/MM2460_g N_VSS_XI39/MM2460_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2443 XI39/NET11098 N_NET256_XI39/MM2443_g N_VSS_XI39/MM2443_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2524 N_NET485_XI39/MM2524_d N_NET387_XI39/MM2524_g N_VSS_XI39/MM2524_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2507 XI39/NET11418 N_NET388_XI39/MM2507_g N_VSS_XI39/MM2507_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2531 N_NET485_XI39/MM2531_d N_NET389_XI39/MM2531_g N_VSS_XI39/MM2531_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2554 XI39/NET11606 N_NET390_XI39/MM2554_g N_VSS_XI39/MM2554_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2211 N_NET485_XI39/MM2211_d N_NET391_XI39/MM2211_g N_VSS_XI39/MM2211_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2234 XI39/NET10418 N_NET262_XI39/MM2234_g N_VSS_XI39/MM2234_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2204 N_NET485_XI39/MM2204_d N_NET263_XI39/MM2204_g N_VSS_XI39/MM2204_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2187 XI39/NET10598 N_NET264_XI39/MM2187_g N_VSS_XI39/MM2187_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2268 N_NET485_XI39/MM2268_d N_NET265_XI39/MM2268_g N_VSS_XI39/MM2268_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2251 XI39/NET10350 N_NET396_XI39/MM2251_g N_VSS_XI39/MM2251_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2275 N_NET485_XI39/MM2275_d N_NET267_XI39/MM2275_g N_VSS_XI39/MM2275_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2298 XI39/NET10170 N_NET268_XI39/MM2298_g N_VSS_XI39/MM2298_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2140 N_NET485_XI39/MM2140_d N_NET269_XI39/MM2140_g N_VSS_XI39/MM2140_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2123 XI39/NET9834 N_NET270_XI39/MM2123_g N_VSS_XI39/MM2123_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2147 N_NET485_XI39/MM2147_d N_NET401_XI39/MM2147_g N_VSS_XI39/MM2147_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2170 XI39/NET9654 N_NET272_XI39/MM2170_g N_VSS_XI39/MM2170_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2083 N_NET485_XI39/MM2083_d N_NET273_XI39/MM2083_g N_VSS_XI39/MM2083_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2106 XI39/NET9906 N_NET404_XI39/MM2106_g N_VSS_XI39/MM2106_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2076 N_NET485_XI39/MM2076_d N_NET405_XI39/MM2076_g N_VSS_XI39/MM2076_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM8 XI39/NET10074 N_NET0390_XI39/MM8_g N_VSS_XI39/MM8_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3414 XI39/NET5566 N_NET0133_XI39/MM3414_g N_VSS_XI39/MM3414_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3394 N_NET486_XI39/MM3394_d N_NET280_XI39/MM3394_g N_VSS_XI39/MM3394_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3429 XI39/NET5506 N_NET281_XI39/MM3429_g N_VSS_XI39/MM3429_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3452 N_NET486_XI39/MM3452_d N_NET282_XI39/MM3452_g N_VSS_XI39/MM3452_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3366 XI39/NET5758 N_NET153_XI39/MM3366_g N_VSS_XI39/MM3366_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3389 N_NET486_XI39/MM3389_d N_NET284_XI39/MM3389_g N_VSS_XI39/MM3389_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3351 XI39/NET3518 N_NET285_XI39/MM3351_g N_VSS_XI39/MM3351_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3330 N_NET486_XI39/MM3330_d N_NET286_XI39/MM3330_g N_VSS_XI39/MM3330_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3493 XI39/NET5250 N_NET287_XI39/MM3493_g N_VSS_XI39/MM3493_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3516 N_NET486_XI39/MM3516_d N_NET158_XI39/MM3516_g N_VSS_XI39/MM3516_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3478 XI39/NET5310 N_NET159_XI39/MM3478_g N_VSS_XI39/MM3478_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3457 N_NET486_XI39/MM3457_d N_NET160_XI39/MM3457_g N_VSS_XI39/MM3457_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3542 XI39/NET5054 N_NET291_XI39/MM3542_g N_VSS_XI39/MM3542_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3521 N_NET486_XI39/MM3521_d N_NET162_XI39/MM3521_g N_VSS_XI39/MM3521_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3557 XI39/NET4994 N_NET293_XI39/MM3557_g N_VSS_XI39/MM3557_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3580 N_NET486_XI39/MM3580_d N_NET294_XI39/MM3580_g N_VSS_XI39/MM3580_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3238 XI39/NET3970 N_NET295_XI39/MM3238_g N_VSS_XI39/MM3238_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3261 N_NET486_XI39/MM3261_d N_NET296_XI39/MM3261_g N_VSS_XI39/MM3261_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3223 XI39/NET4030 N_NET297_XI39/MM3223_g N_VSS_XI39/MM3223_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3202 N_NET486_XI39/MM3202_d N_NET298_XI39/MM3202_g N_VSS_XI39/MM3202_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3287 XI39/NET3774 N_NET299_XI39/MM3287_g N_VSS_XI39/MM3287_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3266 N_NET486_XI39/MM3266_d N_NET170_XI39/MM3266_g N_VSS_XI39/MM3266_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3302 XI39/NET3714 N_NET171_XI39/MM3302_g N_VSS_XI39/MM3302_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3325 N_NET486_XI39/MM3325_d N_NET172_XI39/MM3325_g N_VSS_XI39/MM3325_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3159 XI39/NET4286 N_NET303_XI39/MM3159_g N_VSS_XI39/MM3159_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3138 N_NET486_XI39/MM3138_d N_NET304_XI39/MM3138_g N_VSS_XI39/MM3138_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3174 XI39/NET4226 N_NET305_XI39/MM3174_g N_VSS_XI39/MM3174_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3197 N_NET486_XI39/MM3197_d N_NET306_XI39/MM3197_g N_VSS_XI39/MM3197_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3110 XI39/NET4482 N_NET307_XI39/MM3110_g N_VSS_XI39/MM3110_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3133 N_NET486_XI39/MM3133_d N_NET308_XI39/MM3133_g N_VSS_XI39/MM3133_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3095 XI39/NET4542 N_NET309_XI39/MM3095_g N_VSS_XI39/MM3095_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3074 N_NET486_XI39/MM3074_d N_NET310_XI39/MM3074_g N_VSS_XI39/MM3074_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3839 XI39/NET6166 N_NET311_XI39/MM3839_g N_VSS_XI39/MM3839_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3862 N_NET486_XI39/MM3862_d N_NET312_XI39/MM3862_g N_VSS_XI39/MM3862_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3986 XI39/NET7374 N_NET313_XI39/MM3986_g N_VSS_XI39/MM3986_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3965 N_NET486_XI39/MM3965_d N_NET314_XI39/MM3965_g N_VSS_XI39/MM3965_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3888 XI39/NET5970 N_NET315_XI39/MM3888_g N_VSS_XI39/MM3888_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3867 N_NET486_XI39/MM3867_d N_NET316_XI39/MM3867_g N_VSS_XI39/MM3867_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3903 XI39/NET5910 N_NET317_XI39/MM3903_g N_VSS_XI39/MM3903_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3926 N_NET486_XI39/MM3926_d N_NET318_XI39/MM3926_g N_VSS_XI39/MM3926_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4066 XI39/NET7054 N_NET319_XI39/MM4066_g N_VSS_XI39/MM4066_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4045 N_NET486_XI39/MM4045_d N_NET320_XI39/MM4045_g N_VSS_XI39/MM4045_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3941 XI39/NET7554 N_NET321_XI39/MM3941_g N_VSS_XI39/MM3941_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3960 N_NET486_XI39/MM3960_d N_NET192_XI39/MM3960_g N_VSS_XI39/MM3960_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4017 XI39/NET7250 N_NET193_XI39/MM4017_g N_VSS_XI39/MM4017_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4040 N_NET486_XI39/MM4040_d N_NET194_XI39/MM4040_g N_VSS_XI39/MM4040_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4008 XI39/NET7286 N_NET195_XI39/MM4008_g N_VSS_XI39/MM4008_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4075 N_NET486_XI39/MM4075_d N_NET196_XI39/MM4075_g N_VSS_XI39/MM4075_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3798 XI39/NET6330 N_NET197_XI39/MM3798_g N_VSS_XI39/MM3798_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3777 N_NET486_XI39/MM3777_d N_NET198_XI39/MM3777_g N_VSS_XI39/MM3777_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3813 XI39/NET6270 N_NET199_XI39/MM3813_g N_VSS_XI39/MM3813_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3836 N_NET486_XI39/MM3836_d N_NET200_XI39/MM3836_g N_VSS_XI39/MM3836_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3749 XI39/NET6526 N_NET331_XI39/MM3749_g N_VSS_XI39/MM3749_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3772 N_NET486_XI39/MM3772_d N_NET332_XI39/MM3772_g N_VSS_XI39/MM3772_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3734 XI39/NET6586 N_NET203_XI39/MM3734_g N_VSS_XI39/MM3734_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3713 N_NET486_XI39/MM3713_d N_NET204_XI39/MM3713_g N_VSS_XI39/MM3713_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3621 XI39/NET4738 N_NET205_XI39/MM3621_g N_VSS_XI39/MM3621_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3644 N_NET486_XI39/MM3644_d N_NET206_XI39/MM3644_g N_VSS_XI39/MM3644_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3606 XI39/NET4798 N_NET207_XI39/MM3606_g N_VSS_XI39/MM3606_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3585 N_NET486_XI39/MM3585_d N_NET338_XI39/MM3585_g N_VSS_XI39/MM3585_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3670 XI39/NET6842 N_NET339_XI39/MM3670_g N_VSS_XI39/MM3670_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3649 N_NET486_XI39/MM3649_d N_NET340_XI39/MM3649_g N_VSS_XI39/MM3649_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3686 XI39/NET6778 N_NET211_XI39/MM3686_g N_VSS_XI39/MM3686_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3701 N_NET486_XI39/MM3701_d N_NET212_XI39/MM3701_g N_VSS_XI39/MM3701_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2726 XI39/NET8958 N_NET214_XI39/MM2726_g N_VSS_XI39/MM2726_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2749 N_NET486_XI39/MM2749_d N_NET215_XI39/MM2749_g N_VSS_XI39/MM2749_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2711 XI39/NET9018 N_NET216_XI39/MM2711_g N_VSS_XI39/MM2711_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2690 N_NET486_XI39/MM2690_d N_NET346_XI39/MM2690_g N_VSS_XI39/MM2690_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2775 XI39/NET8766 N_NET347_XI39/MM2775_g N_VSS_XI39/MM2775_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2754 N_NET486_XI39/MM2754_d N_NET348_XI39/MM2754_g N_VSS_XI39/MM2754_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2790 XI39/NET8706 N_NET349_XI39/MM2790_g N_VSS_XI39/MM2790_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2813 N_NET486_XI39/MM2813_d N_NET350_XI39/MM2813_g N_VSS_XI39/MM2813_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2647 XI39/NET9274 N_NET351_XI39/MM2647_g N_VSS_XI39/MM2647_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2626 N_NET486_XI39/MM2626_d N_NET352_XI39/MM2626_g N_VSS_XI39/MM2626_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2662 XI39/NET9214 N_NET224_XI39/MM2662_g N_VSS_XI39/MM2662_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2685 N_NET486_XI39/MM2685_d N_NET225_XI39/MM2685_g N_VSS_XI39/MM2685_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2598 XI39/NET9470 N_NET226_XI39/MM2598_g N_VSS_XI39/MM2598_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2621 N_NET486_XI39/MM2621_d N_NET356_XI39/MM2621_g N_VSS_XI39/MM2621_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2583 XI39/NET9530 N_NET357_XI39/MM2583_g N_VSS_XI39/MM2583_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2562 N_NET486_XI39/MM2562_d N_NET358_XI39/MM2562_g N_VSS_XI39/MM2562_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2903 XI39/NET8254 N_NET230_XI39/MM2903_g N_VSS_XI39/MM2903_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2882 N_NET486_XI39/MM2882_d N_NET360_XI39/MM2882_g N_VSS_XI39/MM2882_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2918 XI39/NET8194 N_NET361_XI39/MM2918_g N_VSS_XI39/MM2918_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2941 N_NET486_XI39/MM2941_d N_NET233_XI39/MM2941_g N_VSS_XI39/MM2941_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2854 XI39/NET8450 N_NET234_XI39/MM2854_g N_VSS_XI39/MM2854_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2877 N_NET486_XI39/MM2877_d N_NET235_XI39/MM2877_g N_VSS_XI39/MM2877_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2839 XI39/NET8510 N_NET365_XI39/MM2839_g N_VSS_XI39/MM2839_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2818 N_NET486_XI39/MM2818_d N_NET366_XI39/MM2818_g N_VSS_XI39/MM2818_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2982 XI39/NET7938 N_NET367_XI39/MM2982_g N_VSS_XI39/MM2982_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3005 N_NET486_XI39/MM3005_d N_NET368_XI39/MM3005_g N_VSS_XI39/MM3005_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2967 XI39/NET7998 N_NET369_XI39/MM2967_g N_VSS_XI39/MM2967_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2946 N_NET486_XI39/MM2946_d N_NET370_XI39/MM2946_g N_VSS_XI39/MM2946_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3031 XI39/NET7742 N_NET371_XI39/MM3031_g N_VSS_XI39/MM3031_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3010 N_NET486_XI39/MM3010_d N_NET242_XI39/MM3010_g N_VSS_XI39/MM3010_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3046 XI39/NET7682 N_NET373_XI39/MM3046_g N_VSS_XI39/MM3046_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3069 N_NET486_XI39/MM3069_d N_NET244_XI39/MM3069_g N_VSS_XI39/MM3069_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2385 XI39/NET10682 N_NET375_XI39/MM2385_g N_VSS_XI39/MM2385_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2370 N_NET486_XI39/MM2370_d N_NET376_XI39/MM2370_g N_VSS_XI39/MM2370_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2406 XI39/NET11246 N_NET377_XI39/MM2406_g N_VSS_XI39/MM2406_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2429 N_NET486_XI39/MM2429_d N_NET378_XI39/MM2429_g N_VSS_XI39/MM2429_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2342 XI39/NET10854 N_NET379_XI39/MM2342_g N_VSS_XI39/MM2342_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2365 N_NET486_XI39/MM2365_d N_NET380_XI39/MM2365_g N_VSS_XI39/MM2365_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2327 XI39/NET10914 N_NET381_XI39/MM2327_g N_VSS_XI39/MM2327_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2306 N_NET486_XI39/MM2306_d N_NET382_XI39/MM2306_g N_VSS_XI39/MM2306_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2472 XI39/NET11558 N_NET383_XI39/MM2472_g N_VSS_XI39/MM2472_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2493 N_NET486_XI39/MM2493_d N_NET384_XI39/MM2493_g N_VSS_XI39/MM2493_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2455 XI39/NET11050 N_NET385_XI39/MM2455_g N_VSS_XI39/MM2455_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2434 N_NET486_XI39/MM2434_d N_NET256_XI39/MM2434_g N_VSS_XI39/MM2434_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2519 XI39/NET11370 N_NET387_XI39/MM2519_g N_VSS_XI39/MM2519_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2498 N_NET486_XI39/MM2498_d N_NET388_XI39/MM2498_g N_VSS_XI39/MM2498_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2528 XI39/NET11334 N_NET389_XI39/MM2528_g N_VSS_XI39/MM2528_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2557 N_NET486_XI39/MM2557_d N_NET390_XI39/MM2557_g N_VSS_XI39/MM2557_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2214 XI39/NET10494 N_NET391_XI39/MM2214_g N_VSS_XI39/MM2214_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2237 N_NET486_XI39/MM2237_d N_NET262_XI39/MM2237_g N_VSS_XI39/MM2237_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2199 XI39/NET10554 N_NET263_XI39/MM2199_g N_VSS_XI39/MM2199_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2178 N_NET486_XI39/MM2178_d N_NET264_XI39/MM2178_g N_VSS_XI39/MM2178_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2263 XI39/NET10306 N_NET265_XI39/MM2263_g N_VSS_XI39/MM2263_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2242 N_NET486_XI39/MM2242_d N_NET396_XI39/MM2242_g N_VSS_XI39/MM2242_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2278 XI39/NET10246 N_NET267_XI39/MM2278_g N_VSS_XI39/MM2278_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2301 N_NET486_XI39/MM2301_d N_NET268_XI39/MM2301_g N_VSS_XI39/MM2301_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2135 XI39/NET9790 N_NET269_XI39/MM2135_g N_VSS_XI39/MM2135_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2114 N_NET486_XI39/MM2114_d N_NET270_XI39/MM2114_g N_VSS_XI39/MM2114_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2150 XI39/NET9730 N_NET401_XI39/MM2150_g N_VSS_XI39/MM2150_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2173 N_NET486_XI39/MM2173_d N_NET272_XI39/MM2173_g N_VSS_XI39/MM2173_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2086 XI39/NET9982 N_NET273_XI39/MM2086_g N_VSS_XI39/MM2086_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2109 N_NET486_XI39/MM2109_d N_NET404_XI39/MM2109_g N_VSS_XI39/MM2109_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2073 XI39/NET10106 N_NET405_XI39/MM2073_g N_VSS_XI39/MM2073_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM13 N_NET486_XI39/MM13_d N_NET0390_XI39/MM13_g N_VSS_XI39/MM13_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI54/XI1/XI10/MM5 N_DOUT<1>_XI54/XI1/XI10/MM5_d
+ N_XI54/XI1/NET9_XI54/XI1/XI10/MM5_g N_VSS_XI54/XI1/XI10/MM5_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=1.68025e-13
+ AS=2.303e-13 PD=7.15e-07 PS=1.45e-06
mXI54/XI1/XI9/MM5 N_XI54/NET16_XI54/XI1/XI9/MM5_d N_DOUT<1>_XI54/XI1/XI9/MM5_g
+ N_VSS_XI54/XI1/XI9/MM5_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.68025e-13 AS=2.303e-13 PD=7.15e-07 PS=1.45e-06
mXI54/XI1/XI10/MM4 N_DOUT<1>_XI54/XI1/XI10/MM4_d
+ N_XI54/NET16_XI54/XI1/XI10/MM4_g N_VSS_XI54/XI1/XI10/MM4_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=1.68025e-13
+ AS=2.3265e-13 PD=7.15e-07 PS=1.46e-06
mXI54/XI1/XI9/MM4 N_XI54/NET16_XI54/XI1/XI9/MM4_d
+ N_XI54/XI1/NET10_XI54/XI1/XI9/MM4_g N_VSS_XI54/XI1/XI9/MM4_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=1.68025e-13
+ AS=2.3265e-13 PD=7.15e-07 PS=1.46e-06
mXI29/XI1/MM45 N_NET487_XI29/XI1/MM45_d N_XI29/XI1/NET219_XI29/XI1/MM45_g
+ N_NET065_XI29/XI1/MM45_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI29/XI1/XI14/MM1 N_XI29/XI1/NET219_XI29/XI1/XI14/MM1_d
+ N_NET464_XI29/XI1/XI14/MM1_g N_VSS_XI29/XI1/XI14/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI29/XI1/MM46 N_NET0395_XI29/XI1/MM46_d N_XI29/XI1/NET207_XI29/XI1/MM46_g
+ N_NET065_XI29/XI1/MM46_s N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI29/XI1/XI15/MM1 N_XI29/XI1/NET207_XI29/XI1/XI15/MM1_d
+ N_NET463_XI29/XI1/XI15/MM1_g N_VSS_XI29/XI1/XI15/MM1_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI39/MM3421 N_NET487_XI39/MM3421_d N_NET0133_XI39/MM3421_g N_VSS_XI39/MM3421_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3405 XI39/NET5602 N_NET280_XI39/MM3405_g N_VSS_XI39/MM3405_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3424 N_NET487_XI39/MM3424_d N_NET281_XI39/MM3424_g N_VSS_XI39/MM3424_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3451 XI39/NET5418 N_NET282_XI39/MM3451_g N_VSS_XI39/MM3451_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3361 N_NET487_XI39/MM3361_d N_NET153_XI39/MM3361_g N_VSS_XI39/MM3361_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3388 XI39/NET5670 N_NET284_XI39/MM3388_g N_VSS_XI39/MM3388_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3358 N_NET487_XI39/MM3358_d N_NET285_XI39/MM3358_g N_VSS_XI39/MM3358_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3329 XI39/NET3606 N_NET286_XI39/MM3329_g N_VSS_XI39/MM3329_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3488 N_NET487_XI39/MM3488_d N_NET287_XI39/MM3488_g N_VSS_XI39/MM3488_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3515 XI39/NET5162 N_NET158_XI39/MM3515_g N_VSS_XI39/MM3515_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3485 N_NET487_XI39/MM3485_d N_NET159_XI39/MM3485_g N_VSS_XI39/MM3485_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3468 XI39/NET5350 N_NET160_XI39/MM3468_g N_VSS_XI39/MM3468_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3549 N_NET487_XI39/MM3549_d N_NET291_XI39/MM3549_g N_VSS_XI39/MM3549_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3532 XI39/NET5094 N_NET162_XI39/MM3532_g N_VSS_XI39/MM3532_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3552 N_NET487_XI39/MM3552_d N_NET293_XI39/MM3552_g N_VSS_XI39/MM3552_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3579 XI39/NET4906 N_NET294_XI39/MM3579_g N_VSS_XI39/MM3579_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3233 N_NET487_XI39/MM3233_d N_NET295_XI39/MM3233_g N_VSS_XI39/MM3233_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3260 XI39/NET3882 N_NET296_XI39/MM3260_g N_VSS_XI39/MM3260_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3230 N_NET487_XI39/MM3230_d N_NET297_XI39/MM3230_g N_VSS_XI39/MM3230_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3213 XI39/NET4070 N_NET298_XI39/MM3213_g N_VSS_XI39/MM3213_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3294 N_NET487_XI39/MM3294_d N_NET299_XI39/MM3294_g N_VSS_XI39/MM3294_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3277 XI39/NET3814 N_NET170_XI39/MM3277_g N_VSS_XI39/MM3277_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3297 N_NET487_XI39/MM3297_d N_NET171_XI39/MM3297_g N_VSS_XI39/MM3297_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3324 XI39/NET3626 N_NET172_XI39/MM3324_g N_VSS_XI39/MM3324_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3166 N_NET487_XI39/MM3166_d N_NET303_XI39/MM3166_g N_VSS_XI39/MM3166_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3149 XI39/NET4326 N_NET304_XI39/MM3149_g N_VSS_XI39/MM3149_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3169 N_NET487_XI39/MM3169_d N_NET305_XI39/MM3169_g N_VSS_XI39/MM3169_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3196 XI39/NET4138 N_NET306_XI39/MM3196_g N_VSS_XI39/MM3196_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3105 N_NET487_XI39/MM3105_d N_NET307_XI39/MM3105_g N_VSS_XI39/MM3105_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3132 XI39/NET4394 N_NET308_XI39/MM3132_g N_VSS_XI39/MM3132_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3102 N_NET487_XI39/MM3102_d N_NET309_XI39/MM3102_g N_VSS_XI39/MM3102_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3085 XI39/NET4582 N_NET310_XI39/MM3085_g N_VSS_XI39/MM3085_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3996 N_NET487_XI39/MM3996_d N_NET311_XI39/MM3996_g N_VSS_XI39/MM3996_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3861 XI39/NET6078 N_NET312_XI39/MM3861_g N_VSS_XI39/MM3861_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3993 N_NET487_XI39/MM3993_d N_NET313_XI39/MM3993_g N_VSS_XI39/MM3993_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3976 XI39/NET7414 N_NET314_XI39/MM3976_g N_VSS_XI39/MM3976_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3895 N_NET487_XI39/MM3895_d N_NET315_XI39/MM3895_g N_VSS_XI39/MM3895_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3878 XI39/NET6010 N_NET316_XI39/MM3878_g N_VSS_XI39/MM3878_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3898 N_NET487_XI39/MM3898_d N_NET317_XI39/MM3898_g N_VSS_XI39/MM3898_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3925 XI39/NET5822 N_NET318_XI39/MM3925_g N_VSS_XI39/MM3925_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3929 N_NET487_XI39/MM3929_d N_NET319_XI39/MM3929_g N_VSS_XI39/MM3929_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4056 XI39/NET7094 N_NET320_XI39/MM4056_g N_VSS_XI39/MM4056_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3932 N_NET487_XI39/MM3932_d N_NET321_XI39/MM3932_g N_VSS_XI39/MM3932_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3959 XI39/NET7482 N_NET192_XI39/MM3959_g N_VSS_XI39/MM3959_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4012 N_NET487_XI39/MM4012_d N_NET193_XI39/MM4012_g N_VSS_XI39/MM4012_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4039 XI39/NET7162 N_NET194_XI39/MM4039_g N_VSS_XI39/MM4039_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4009 N_NET487_XI39/MM4009_d N_NET195_XI39/MM4009_g N_VSS_XI39/MM4009_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4086 XI39/NET6974 N_NET196_XI39/MM4086_g N_VSS_XI39/MM4086_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3805 N_NET487_XI39/MM3805_d N_NET197_XI39/MM3805_g N_VSS_XI39/MM3805_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3788 XI39/NET6370 N_NET198_XI39/MM3788_g N_VSS_XI39/MM3788_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3808 N_NET487_XI39/MM3808_d N_NET199_XI39/MM3808_g N_VSS_XI39/MM3808_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3835 XI39/NET6182 N_NET200_XI39/MM3835_g N_VSS_XI39/MM3835_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3744 N_NET487_XI39/MM3744_d N_NET331_XI39/MM3744_g N_VSS_XI39/MM3744_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3771 XI39/NET6438 N_NET332_XI39/MM3771_g N_VSS_XI39/MM3771_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3741 N_NET487_XI39/MM3741_d N_NET203_XI39/MM3741_g N_VSS_XI39/MM3741_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3724 XI39/NET6626 N_NET204_XI39/MM3724_g N_VSS_XI39/MM3724_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3616 N_NET487_XI39/MM3616_d N_NET205_XI39/MM3616_g N_VSS_XI39/MM3616_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3643 XI39/NET4650 N_NET206_XI39/MM3643_g N_VSS_XI39/MM3643_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3613 N_NET487_XI39/MM3613_d N_NET207_XI39/MM3613_g N_VSS_XI39/MM3613_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3596 XI39/NET4838 N_NET338_XI39/MM3596_g N_VSS_XI39/MM3596_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3677 N_NET487_XI39/MM3677_d N_NET339_XI39/MM3677_g N_VSS_XI39/MM3677_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3660 XI39/NET6882 N_NET340_XI39/MM3660_g N_VSS_XI39/MM3660_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3709 N_NET487_XI39/MM3709_d N_NET211_XI39/MM3709_g N_VSS_XI39/MM3709_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3700 XI39/NET6722 N_NET212_XI39/MM3700_g N_VSS_XI39/MM3700_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2721 N_NET487_XI39/MM2721_d N_NET214_XI39/MM2721_g N_VSS_XI39/MM2721_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2748 XI39/NET8874 N_NET215_XI39/MM2748_g N_VSS_XI39/MM2748_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2718 N_NET487_XI39/MM2718_d N_NET216_XI39/MM2718_g N_VSS_XI39/MM2718_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2701 XI39/NET9058 N_NET346_XI39/MM2701_g N_VSS_XI39/MM2701_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2782 N_NET487_XI39/MM2782_d N_NET347_XI39/MM2782_g N_VSS_XI39/MM2782_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2765 XI39/NET8806 N_NET348_XI39/MM2765_g N_VSS_XI39/MM2765_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2785 N_NET487_XI39/MM2785_d N_NET349_XI39/MM2785_g N_VSS_XI39/MM2785_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2812 XI39/NET8618 N_NET350_XI39/MM2812_g N_VSS_XI39/MM2812_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2654 N_NET487_XI39/MM2654_d N_NET351_XI39/MM2654_g N_VSS_XI39/MM2654_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2637 XI39/NET9314 N_NET352_XI39/MM2637_g N_VSS_XI39/MM2637_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2657 N_NET487_XI39/MM2657_d N_NET224_XI39/MM2657_g N_VSS_XI39/MM2657_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2684 XI39/NET9126 N_NET225_XI39/MM2684_g N_VSS_XI39/MM2684_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2593 N_NET487_XI39/MM2593_d N_NET226_XI39/MM2593_g N_VSS_XI39/MM2593_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2620 XI39/NET9382 N_NET356_XI39/MM2620_g N_VSS_XI39/MM2620_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2590 N_NET487_XI39/MM2590_d N_NET357_XI39/MM2590_g N_VSS_XI39/MM2590_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2573 XI39/NET9570 N_NET358_XI39/MM2573_g N_VSS_XI39/MM2573_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2910 N_NET487_XI39/MM2910_d N_NET230_XI39/MM2910_g N_VSS_XI39/MM2910_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2893 XI39/NET8294 N_NET360_XI39/MM2893_g N_VSS_XI39/MM2893_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2913 N_NET487_XI39/MM2913_d N_NET361_XI39/MM2913_g N_VSS_XI39/MM2913_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2940 XI39/NET8106 N_NET233_XI39/MM2940_g N_VSS_XI39/MM2940_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2849 N_NET487_XI39/MM2849_d N_NET234_XI39/MM2849_g N_VSS_XI39/MM2849_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2876 XI39/NET8362 N_NET235_XI39/MM2876_g N_VSS_XI39/MM2876_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2846 N_NET487_XI39/MM2846_d N_NET365_XI39/MM2846_g N_VSS_XI39/MM2846_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2829 XI39/NET8550 N_NET366_XI39/MM2829_g N_VSS_XI39/MM2829_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2977 N_NET487_XI39/MM2977_d N_NET367_XI39/MM2977_g N_VSS_XI39/MM2977_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3004 XI39/NET7850 N_NET368_XI39/MM3004_g N_VSS_XI39/MM3004_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2974 N_NET487_XI39/MM2974_d N_NET369_XI39/MM2974_g N_VSS_XI39/MM2974_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2957 XI39/NET8038 N_NET370_XI39/MM2957_g N_VSS_XI39/MM2957_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3038 N_NET487_XI39/MM3038_d N_NET371_XI39/MM3038_g N_VSS_XI39/MM3038_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3021 XI39/NET7782 N_NET242_XI39/MM3021_g N_VSS_XI39/MM3021_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3041 N_NET487_XI39/MM3041_d N_NET373_XI39/MM3041_g N_VSS_XI39/MM3041_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3068 XI39/NET7594 N_NET244_XI39/MM3068_g N_VSS_XI39/MM3068_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2398 N_NET487_XI39/MM2398_d N_NET375_XI39/MM2398_g N_VSS_XI39/MM2398_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2381 XI39/NET10698 N_NET376_XI39/MM2381_g N_VSS_XI39/MM2381_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2401 N_NET487_XI39/MM2401_d N_NET377_XI39/MM2401_g N_VSS_XI39/MM2401_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2428 XI39/NET11158 N_NET378_XI39/MM2428_g N_VSS_XI39/MM2428_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2337 N_NET487_XI39/MM2337_d N_NET379_XI39/MM2337_g N_VSS_XI39/MM2337_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2364 XI39/NET10766 N_NET380_XI39/MM2364_g N_VSS_XI39/MM2364_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2334 N_NET487_XI39/MM2334_d N_NET381_XI39/MM2334_g N_VSS_XI39/MM2334_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2317 XI39/NET10954 N_NET382_XI39/MM2317_g N_VSS_XI39/MM2317_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2465 N_NET487_XI39/MM2465_d N_NET383_XI39/MM2465_g N_VSS_XI39/MM2465_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2492 XI39/NET11478 N_NET384_XI39/MM2492_g N_VSS_XI39/MM2492_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2462 N_NET487_XI39/MM2462_d N_NET385_XI39/MM2462_g N_VSS_XI39/MM2462_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2445 XI39/NET11090 N_NET256_XI39/MM2445_g N_VSS_XI39/MM2445_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2526 N_NET487_XI39/MM2526_d N_NET387_XI39/MM2526_g N_VSS_XI39/MM2526_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2509 XI39/NET11410 N_NET388_XI39/MM2509_g N_VSS_XI39/MM2509_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2529 N_NET487_XI39/MM2529_d N_NET389_XI39/MM2529_g N_VSS_XI39/MM2529_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2556 XI39/NET11598 N_NET390_XI39/MM2556_g N_VSS_XI39/MM2556_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2209 N_NET487_XI39/MM2209_d N_NET391_XI39/MM2209_g N_VSS_XI39/MM2209_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2236 XI39/NET10410 N_NET262_XI39/MM2236_g N_VSS_XI39/MM2236_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2206 N_NET487_XI39/MM2206_d N_NET263_XI39/MM2206_g N_VSS_XI39/MM2206_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2189 XI39/NET10590 N_NET264_XI39/MM2189_g N_VSS_XI39/MM2189_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2270 N_NET487_XI39/MM2270_d N_NET265_XI39/MM2270_g N_VSS_XI39/MM2270_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2253 XI39/NET10342 N_NET396_XI39/MM2253_g N_VSS_XI39/MM2253_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2273 N_NET487_XI39/MM2273_d N_NET267_XI39/MM2273_g N_VSS_XI39/MM2273_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2300 XI39/NET10162 N_NET268_XI39/MM2300_g N_VSS_XI39/MM2300_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2142 N_NET487_XI39/MM2142_d N_NET269_XI39/MM2142_g N_VSS_XI39/MM2142_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2125 XI39/NET9826 N_NET270_XI39/MM2125_g N_VSS_XI39/MM2125_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2145 N_NET487_XI39/MM2145_d N_NET401_XI39/MM2145_g N_VSS_XI39/MM2145_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2172 XI39/NET9646 N_NET272_XI39/MM2172_g N_VSS_XI39/MM2172_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2081 N_NET487_XI39/MM2081_d N_NET273_XI39/MM2081_g N_VSS_XI39/MM2081_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2108 XI39/NET9898 N_NET404_XI39/MM2108_g N_VSS_XI39/MM2108_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2078 N_NET487_XI39/MM2078_d N_NET405_XI39/MM2078_g N_VSS_XI39/MM2078_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM0 XI39/NET10042 N_NET0390_XI39/MM0_g N_VSS_XI39/MM0_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3422 XI39/NET5534 N_NET0133_XI39/MM3422_g N_VSS_XI39/MM3422_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3392 N_NET0395_XI39/MM3392_d N_NET280_XI39/MM3392_g N_VSS_XI39/MM3392_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3437 XI39/NET5474 N_NET281_XI39/MM3437_g N_VSS_XI39/MM3437_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3454 N_NET0395_XI39/MM3454_d N_NET282_XI39/MM3454_g N_VSS_XI39/MM3454_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3374 XI39/NET5726 N_NET153_XI39/MM3374_g N_VSS_XI39/MM3374_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3391 N_NET0395_XI39/MM3391_d N_NET284_XI39/MM3391_g N_VSS_XI39/MM3391_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3359 XI39/NET3486 N_NET285_XI39/MM3359_g N_VSS_XI39/MM3359_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3328 N_NET0395_XI39/MM3328_d N_NET286_XI39/MM3328_g N_VSS_XI39/MM3328_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3501 XI39/NET5218 N_NET287_XI39/MM3501_g N_VSS_XI39/MM3501_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3518 N_NET0395_XI39/MM3518_d N_NET158_XI39/MM3518_g N_VSS_XI39/MM3518_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3486 XI39/NET5278 N_NET159_XI39/MM3486_g N_VSS_XI39/MM3486_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3455 N_NET0395_XI39/MM3455_d N_NET160_XI39/MM3455_g N_VSS_XI39/MM3455_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3550 XI39/NET5022 N_NET291_XI39/MM3550_g N_VSS_XI39/MM3550_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3519 N_NET0395_XI39/MM3519_d N_NET162_XI39/MM3519_g N_VSS_XI39/MM3519_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3565 XI39/NET4962 N_NET293_XI39/MM3565_g N_VSS_XI39/MM3565_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3582 N_NET0395_XI39/MM3582_d N_NET294_XI39/MM3582_g N_VSS_XI39/MM3582_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3246 XI39/NET3938 N_NET295_XI39/MM3246_g N_VSS_XI39/MM3246_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3263 N_NET0395_XI39/MM3263_d N_NET296_XI39/MM3263_g N_VSS_XI39/MM3263_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3231 XI39/NET3998 N_NET297_XI39/MM3231_g N_VSS_XI39/MM3231_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3200 N_NET0395_XI39/MM3200_d N_NET298_XI39/MM3200_g N_VSS_XI39/MM3200_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3295 XI39/NET3742 N_NET299_XI39/MM3295_g N_VSS_XI39/MM3295_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3264 N_NET0395_XI39/MM3264_d N_NET170_XI39/MM3264_g N_VSS_XI39/MM3264_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3310 XI39/NET3682 N_NET171_XI39/MM3310_g N_VSS_XI39/MM3310_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3327 N_NET0395_XI39/MM3327_d N_NET172_XI39/MM3327_g N_VSS_XI39/MM3327_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3167 XI39/NET4254 N_NET303_XI39/MM3167_g N_VSS_XI39/MM3167_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3136 N_NET0395_XI39/MM3136_d N_NET304_XI39/MM3136_g N_VSS_XI39/MM3136_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3182 XI39/NET4194 N_NET305_XI39/MM3182_g N_VSS_XI39/MM3182_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3199 N_NET0395_XI39/MM3199_d N_NET306_XI39/MM3199_g N_VSS_XI39/MM3199_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3118 XI39/NET4450 N_NET307_XI39/MM3118_g N_VSS_XI39/MM3118_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3135 N_NET0395_XI39/MM3135_d N_NET308_XI39/MM3135_g N_VSS_XI39/MM3135_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3103 XI39/NET4510 N_NET309_XI39/MM3103_g N_VSS_XI39/MM3103_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3072 N_NET0395_XI39/MM3072_d N_NET310_XI39/MM3072_g N_VSS_XI39/MM3072_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3847 XI39/NET6134 N_NET311_XI39/MM3847_g N_VSS_XI39/MM3847_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3864 N_NET0395_XI39/MM3864_d N_NET312_XI39/MM3864_g N_VSS_XI39/MM3864_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3994 XI39/NET7342 N_NET313_XI39/MM3994_g N_VSS_XI39/MM3994_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3963 N_NET0395_XI39/MM3963_d N_NET314_XI39/MM3963_g N_VSS_XI39/MM3963_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3896 XI39/NET5938 N_NET315_XI39/MM3896_g N_VSS_XI39/MM3896_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3865 N_NET0395_XI39/MM3865_d N_NET316_XI39/MM3865_g N_VSS_XI39/MM3865_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3911 XI39/NET5878 N_NET317_XI39/MM3911_g N_VSS_XI39/MM3911_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3928 N_NET0395_XI39/MM3928_d N_NET318_XI39/MM3928_g N_VSS_XI39/MM3928_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3930 XI39/NET5802 N_NET319_XI39/MM3930_g N_VSS_XI39/MM3930_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4043 N_NET0395_XI39/MM4043_d N_NET320_XI39/MM4043_g N_VSS_XI39/MM4043_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3933 XI39/NET5790 N_NET321_XI39/MM3933_g N_VSS_XI39/MM3933_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3962 N_NET0395_XI39/MM3962_d N_NET192_XI39/MM3962_g N_VSS_XI39/MM3962_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4025 XI39/NET7218 N_NET193_XI39/MM4025_g N_VSS_XI39/MM4025_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4042 N_NET0395_XI39/MM4042_d N_NET194_XI39/MM4042_g N_VSS_XI39/MM4042_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4094 XI39/NET6942 N_NET195_XI39/MM4094_g N_VSS_XI39/MM4094_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM4073 N_NET0395_XI39/MM4073_d N_NET196_XI39/MM4073_g N_VSS_XI39/MM4073_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3806 XI39/NET6298 N_NET197_XI39/MM3806_g N_VSS_XI39/MM3806_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3775 N_NET0395_XI39/MM3775_d N_NET198_XI39/MM3775_g N_VSS_XI39/MM3775_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3821 XI39/NET6238 N_NET199_XI39/MM3821_g N_VSS_XI39/MM3821_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3838 N_NET0395_XI39/MM3838_d N_NET200_XI39/MM3838_g N_VSS_XI39/MM3838_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3757 XI39/NET6494 N_NET331_XI39/MM3757_g N_VSS_XI39/MM3757_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3774 N_NET0395_XI39/MM3774_d N_NET332_XI39/MM3774_g N_VSS_XI39/MM3774_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3742 XI39/NET6554 N_NET203_XI39/MM3742_g N_VSS_XI39/MM3742_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3711 N_NET0395_XI39/MM3711_d N_NET204_XI39/MM3711_g N_VSS_XI39/MM3711_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3629 XI39/NET4706 N_NET205_XI39/MM3629_g N_VSS_XI39/MM3629_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3646 N_NET0395_XI39/MM3646_d N_NET206_XI39/MM3646_g N_VSS_XI39/MM3646_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3614 XI39/NET4766 N_NET207_XI39/MM3614_g N_VSS_XI39/MM3614_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3583 N_NET0395_XI39/MM3583_d N_NET338_XI39/MM3583_g N_VSS_XI39/MM3583_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3678 XI39/NET6810 N_NET339_XI39/MM3678_g N_VSS_XI39/MM3678_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3647 N_NET0395_XI39/MM3647_d N_NET340_XI39/MM3647_g N_VSS_XI39/MM3647_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3710 XI39/NET6682 N_NET211_XI39/MM3710_g N_VSS_XI39/MM3710_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3703 N_NET0395_XI39/MM3703_d N_NET212_XI39/MM3703_g N_VSS_XI39/MM3703_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2734 XI39/NET8926 N_NET214_XI39/MM2734_g N_VSS_XI39/MM2734_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2751 N_NET0395_XI39/MM2751_d N_NET215_XI39/MM2751_g N_VSS_XI39/MM2751_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2719 XI39/NET8986 N_NET216_XI39/MM2719_g N_VSS_XI39/MM2719_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2688 N_NET0395_XI39/MM2688_d N_NET346_XI39/MM2688_g N_VSS_XI39/MM2688_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2783 XI39/NET8734 N_NET347_XI39/MM2783_g N_VSS_XI39/MM2783_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2752 N_NET0395_XI39/MM2752_d N_NET348_XI39/MM2752_g N_VSS_XI39/MM2752_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2798 XI39/NET8674 N_NET349_XI39/MM2798_g N_VSS_XI39/MM2798_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2815 N_NET0395_XI39/MM2815_d N_NET350_XI39/MM2815_g N_VSS_XI39/MM2815_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2655 XI39/NET9242 N_NET351_XI39/MM2655_g N_VSS_XI39/MM2655_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2624 N_NET0395_XI39/MM2624_d N_NET352_XI39/MM2624_g N_VSS_XI39/MM2624_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2670 XI39/NET9182 N_NET224_XI39/MM2670_g N_VSS_XI39/MM2670_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2687 N_NET0395_XI39/MM2687_d N_NET225_XI39/MM2687_g N_VSS_XI39/MM2687_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2606 XI39/NET9438 N_NET226_XI39/MM2606_g N_VSS_XI39/MM2606_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2623 N_NET0395_XI39/MM2623_d N_NET356_XI39/MM2623_g N_VSS_XI39/MM2623_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2591 XI39/NET9498 N_NET357_XI39/MM2591_g N_VSS_XI39/MM2591_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2560 N_NET0395_XI39/MM2560_d N_NET358_XI39/MM2560_g N_VSS_XI39/MM2560_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2911 XI39/NET8222 N_NET230_XI39/MM2911_g N_VSS_XI39/MM2911_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2880 N_NET0395_XI39/MM2880_d N_NET360_XI39/MM2880_g N_VSS_XI39/MM2880_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2926 XI39/NET8162 N_NET361_XI39/MM2926_g N_VSS_XI39/MM2926_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2943 N_NET0395_XI39/MM2943_d N_NET233_XI39/MM2943_g N_VSS_XI39/MM2943_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2862 XI39/NET8418 N_NET234_XI39/MM2862_g N_VSS_XI39/MM2862_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2879 N_NET0395_XI39/MM2879_d N_NET235_XI39/MM2879_g N_VSS_XI39/MM2879_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2847 XI39/NET8478 N_NET365_XI39/MM2847_g N_VSS_XI39/MM2847_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2816 N_NET0395_XI39/MM2816_d N_NET366_XI39/MM2816_g N_VSS_XI39/MM2816_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2990 XI39/NET7906 N_NET367_XI39/MM2990_g N_VSS_XI39/MM2990_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3007 N_NET0395_XI39/MM3007_d N_NET368_XI39/MM3007_g N_VSS_XI39/MM3007_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2975 XI39/NET7966 N_NET369_XI39/MM2975_g N_VSS_XI39/MM2975_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2944 N_NET0395_XI39/MM2944_d N_NET370_XI39/MM2944_g N_VSS_XI39/MM2944_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3039 XI39/NET7710 N_NET371_XI39/MM3039_g N_VSS_XI39/MM3039_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3008 N_NET0395_XI39/MM3008_d N_NET242_XI39/MM3008_g N_VSS_XI39/MM3008_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3054 XI39/NET7650 N_NET373_XI39/MM3054_g N_VSS_XI39/MM3054_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM3071 N_NET0395_XI39/MM3071_d N_NET244_XI39/MM3071_g N_VSS_XI39/MM3071_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2393 XI39/NET10650 N_NET375_XI39/MM2393_g N_VSS_XI39/MM2393_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2368 N_NET0395_XI39/MM2368_d N_NET376_XI39/MM2368_g N_VSS_XI39/MM2368_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2414 XI39/NET11214 N_NET377_XI39/MM2414_g N_VSS_XI39/MM2414_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2431 N_NET0395_XI39/MM2431_d N_NET378_XI39/MM2431_g N_VSS_XI39/MM2431_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2350 XI39/NET10822 N_NET379_XI39/MM2350_g N_VSS_XI39/MM2350_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2367 N_NET0395_XI39/MM2367_d N_NET380_XI39/MM2367_g N_VSS_XI39/MM2367_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2335 XI39/NET10882 N_NET381_XI39/MM2335_g N_VSS_XI39/MM2335_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2304 N_NET0395_XI39/MM2304_d N_NET382_XI39/MM2304_g N_VSS_XI39/MM2304_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2464 XI39/NET11014 N_NET383_XI39/MM2464_g N_VSS_XI39/MM2464_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2495 N_NET0395_XI39/MM2495_d N_NET384_XI39/MM2495_g N_VSS_XI39/MM2495_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2463 XI39/NET11018 N_NET385_XI39/MM2463_g N_VSS_XI39/MM2463_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2432 N_NET0395_XI39/MM2432_d N_NET256_XI39/MM2432_g N_VSS_XI39/MM2432_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2527 XI39/NET11338 N_NET387_XI39/MM2527_g N_VSS_XI39/MM2527_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2496 N_NET0395_XI39/MM2496_d N_NET388_XI39/MM2496_g N_VSS_XI39/MM2496_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2536 XI39/NET11302 N_NET389_XI39/MM2536_g N_VSS_XI39/MM2536_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2559 N_NET0395_XI39/MM2559_d N_NET390_XI39/MM2559_g N_VSS_XI39/MM2559_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2222 XI39/NET10462 N_NET391_XI39/MM2222_g N_VSS_XI39/MM2222_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2239 N_NET0395_XI39/MM2239_d N_NET262_XI39/MM2239_g N_VSS_XI39/MM2239_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2207 XI39/NET10522 N_NET263_XI39/MM2207_g N_VSS_XI39/MM2207_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2176 N_NET0395_XI39/MM2176_d N_NET264_XI39/MM2176_g N_VSS_XI39/MM2176_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2271 XI39/NET10274 N_NET265_XI39/MM2271_g N_VSS_XI39/MM2271_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2240 N_NET0395_XI39/MM2240_d N_NET396_XI39/MM2240_g N_VSS_XI39/MM2240_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2286 XI39/NET10214 N_NET267_XI39/MM2286_g N_VSS_XI39/MM2286_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2303 N_NET0395_XI39/MM2303_d N_NET268_XI39/MM2303_g N_VSS_XI39/MM2303_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2143 XI39/NET9758 N_NET269_XI39/MM2143_g N_VSS_XI39/MM2143_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2112 N_NET0395_XI39/MM2112_d N_NET270_XI39/MM2112_g N_VSS_XI39/MM2112_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2158 XI39/NET9698 N_NET401_XI39/MM2158_g N_VSS_XI39/MM2158_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2175 N_NET0395_XI39/MM2175_d N_NET272_XI39/MM2175_g N_VSS_XI39/MM2175_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2094 XI39/NET9950 N_NET273_XI39/MM2094_g N_VSS_XI39/MM2094_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2111 N_NET0395_XI39/MM2111_d N_NET404_XI39/MM2111_g N_VSS_XI39/MM2111_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM2065 XI39/NET10010 N_NET405_XI39/MM2065_g N_VSS_XI39/MM2065_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI39/MM15 N_NET0395_XI39/MM15_d N_NET0390_XI39/MM15_g N_VSS_XI39/MM15_s
+ N_VSS_XI42/XI519/XI72/XI21/MM5_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI42/XI519/XI72/XI21/MM6
+ N_XI42/XI519/XI72/XI21/NET21_XI42/XI519/XI72/XI21/MM6_d
+ N_NET127_XI42/XI519/XI72/XI21/MM6_g N_VDD_XI42/XI519/XI72/XI21/MM6_s
+ N_VDD_XI42/XI519/XI72/XI21/MM6_b P_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13
+ AS=2.632e-13 PD=7.2e-07 PS=1.59e-06
mXI42/XI519/XI73/XI21/MM6
+ N_XI42/XI519/XI73/XI21/NET21_XI42/XI519/XI73/XI21/MM6_d
+ N_NET141_XI42/XI519/XI73/XI21/MM6_g N_VDD_XI42/XI519/XI73/XI21/MM6_s
+ N_VDD_XI42/XI519/XI73/XI21/MM6_b P_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13
+ AS=2.632e-13 PD=7.2e-07 PS=1.59e-06
mXI48/XI66/MM0 N_XI48/XI66/NET52_XI48/XI66/MM0_d N_CLK_XI48/XI66/MM0_g
+ N_A<9>_XI48/XI66/MM0_s N_VDD_XI48/XI66/MM0_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI48/XI66/MM1 N_XI48/XI66/NET48_XI48/XI66/MM1_d N_NET90_XI48/XI66/MM1_g
+ N_XI48/XI66/NET52_XI48/XI66/MM1_s N_VDD_XI48/XI66/MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI48/XI65/MM0 N_XI48/XI65/NET52_XI48/XI65/MM0_d N_CLK_XI48/XI65/MM0_g
+ N_A<8>_XI48/XI65/MM0_s N_VDD_XI48/XI66/MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI48/XI65/MM1 N_XI48/XI65/NET48_XI48/XI65/MM1_d N_NET90_XI48/XI65/MM1_g
+ N_XI48/XI65/NET52_XI48/XI65/MM1_s N_VDD_XI48/XI65/MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI48/XI64/MM0 N_XI48/XI64/NET52_XI48/XI64/MM0_d N_CLK_XI48/XI64/MM0_g
+ N_A<7>_XI48/XI64/MM0_s N_VDD_XI48/XI65/MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI48/XI64/MM1 N_XI48/XI64/NET48_XI48/XI64/MM1_d N_NET90_XI48/XI64/MM1_g
+ N_XI48/XI64/NET52_XI48/XI64/MM1_s N_VDD_XI48/XI64/MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI48/XI74/XI3/MM0 N_NET136_XI48/XI74/XI3/MM0_d N_NET135_XI48/XI74/XI3/MM0_g
+ N_VDD_XI48/XI74/XI3/MM0_s N_VDD_XI48/XI66/MM1_b P_18 L=1.8e-07 W=1.85e-06
+ AD=9.435e-13 AS=9.435e-13 PD=2.87e-06 PS=2.87e-06
mXI48/XI73/XI3/MM0 N_NET138_XI48/XI73/XI3/MM0_d N_NET137_XI48/XI73/XI3/MM0_g
+ N_VDD_XI48/XI73/XI3/MM0_s N_VDD_XI48/XI65/MM1_b P_18 L=1.8e-07 W=1.85e-06
+ AD=9.435e-13 AS=9.435e-13 PD=2.87e-06 PS=2.87e-06
mXI48/XI72/XI3/MM0 N_NET140_XI48/XI72/XI3/MM0_d N_NET139_XI48/XI72/XI3/MM0_g
+ N_VDD_XI48/XI72/XI3/MM0_s N_VDD_XI48/XI64/MM1_b P_18 L=1.8e-07 W=1.85e-06
+ AD=9.435e-13 AS=9.435e-13 PD=2.87e-06 PS=2.87e-06
mXI48/XI60/MM1 N_XI48/XI60/NET48_XI48/XI60/MM1_d N_NET90_XI48/XI60/MM1_g
+ N_XI48/XI60/NET52_XI48/XI60/MM1_s N_VDD_XI48/XI60/MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI48/XI60/MM0 N_XI48/XI60/NET52_XI48/XI60/MM0_d N_CLK_XI48/XI60/MM0_g
+ N_A<3>_XI48/XI60/MM0_s N_VDD_XI48/XI60/MM0_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI48/XI61/MM0 N_XI48/XI61/NET52_XI48/XI61/MM0_d N_CLK_XI48/XI61/MM0_g
+ N_A<4>_XI48/XI61/MM0_s N_VDD_XI42/XI519/XI72/XI21/MM6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI48/XI61/MM1 N_XI48/XI61/NET48_XI48/XI61/MM1_d N_NET90_XI48/XI61/MM1_g
+ N_XI48/XI61/NET52_XI48/XI61/MM1_s N_VDD_XI48/XI61/MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI48/XI62/MM1 N_XI48/XI62/NET48_XI48/XI62/MM1_d N_NET90_XI48/XI62/MM1_g
+ N_XI48/XI62/NET52_XI48/XI62/MM1_s N_VDD_XI48/XI62/MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI48/XI62/MM0 N_XI48/XI62/NET52_XI48/XI62/MM0_d N_CLK_XI48/XI62/MM0_g
+ N_A<5>_XI48/XI62/MM0_s N_VDD_XI48/XI62/MM0_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI48/XI63/MM0 N_XI48/XI63/NET52_XI48/XI63/MM0_d N_CLK_XI48/XI63/MM0_g
+ N_A<6>_XI48/XI63/MM0_s N_VDD_XI42/XI519/XI73/XI21/MM6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI48/XI63/MM1 N_XI48/XI63/NET48_XI48/XI63/MM1_d N_NET90_XI48/XI63/MM1_g
+ N_XI48/XI63/NET52_XI48/XI63/MM1_s N_VDD_XI48/XI63/MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI32/XI9/MM0 N_XI32/XI9/NET52_XI32/XI9/MM0_d N_CLK_XI32/XI9/MM0_g
+ N_A<2>_XI32/XI9/MM0_s N_VDD_XI48/XI63/MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI32/XI9/MM1 N_XI32/XI9/NET48_XI32/XI9/MM1_d N_NET90_XI32/XI9/MM1_g
+ N_XI32/XI9/NET52_XI32/XI9/MM1_s N_VDD_XI32/XI9/MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI32/XI8/MM0 N_XI32/XI8/NET52_XI32/XI8/MM0_d N_CLK_XI32/XI8/MM0_g
+ N_A<1>_XI32/XI8/MM0_s N_VDD_XI32/XI9/MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI32/XI8/MM1 N_XI32/XI8/NET48_XI32/XI8/MM1_d N_NET90_XI32/XI8/MM1_g
+ N_XI32/XI8/NET52_XI32/XI8/MM1_s N_VDD_XI32/XI8/MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI32/XI7/MM0 N_XI32/XI7/NET52_XI32/XI7/MM0_d N_CLK_XI32/XI7/MM0_g
+ N_A<0>_XI32/XI7/MM0_s N_VDD_XI32/XI8/MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI32/XI7/MM1 N_XI32/XI7/NET48_XI32/XI7/MM1_d N_NET90_XI32/XI7/MM1_g
+ N_XI32/XI7/NET52_XI32/XI7/MM1_s N_VDD_XI32/XI7/MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI42/XI519/XI72/XI21/MM7 N_XI42/XI519/NET114_XI42/XI519/XI72/XI21/MM7_d
+ N_NET129_XI42/XI519/XI72/XI21/MM7_g
+ N_XI42/XI519/XI72/XI21/NET21_XI42/XI519/XI72/XI21/MM7_s
+ N_VDD_XI42/XI519/XI72/XI21/MM6_b P_18 L=1.8e-07 W=4.7e-07 AD=2.397e-13
+ AS=1.692e-13 PD=1.49e-06 PS=7.2e-07
mXI42/XI519/XI73/XI21/MM7 N_XI42/XI519/NET36_XI42/XI519/XI73/XI21/MM7_d
+ N_NET143_XI42/XI519/XI73/XI21/MM7_g
+ N_XI42/XI519/XI73/XI21/NET21_XI42/XI519/XI73/XI21/MM7_s
+ N_VDD_XI42/XI519/XI73/XI21/MM6_b P_18 L=1.8e-07 W=4.7e-07 AD=2.397e-13
+ AS=1.692e-13 PD=1.49e-06 PS=7.2e-07
mXI56/MM0 N_NET90_XI56/MM0_d N_CLK_XI56/MM0_g N_VDD_XI56/MM0_s
+ N_VDD_XI32/XI7/MM1_b P_18 L=1.8e-07 W=1.85e-06 AD=9.065e-13 AS=9.065e-13
+ PD=2.83e-06 PS=2.83e-06
mXI58/XI164/XI0/MM0 N_XI58/XI164/NET10_XI58/XI164/XI0/MM0_d
+ N_CLK_XI58/XI164/XI0/MM0_g N_VDD_XI58/XI164/XI0/MM0_s N_VDD_XI32/XI7/MM1_b
+ P_18 L=1.8e-07 W=1.85e-06 AD=4.7175e-13 AS=9.065e-13 PD=5.1e-07 PS=2.83e-06
mXI58/XI164/XI0/MM0@2 N_XI58/XI164/NET10_XI58/XI164/XI0/MM0@2_d
+ N_CLK_XI58/XI164/XI0/MM0@2_g N_VDD_XI58/XI164/XI0/MM0@2_s N_VDD_XI32/XI7/MM1_b
+ P_18 L=1.8e-07 W=1.85e-06 AD=4.7175e-13 AS=9.065e-13 PD=5.1e-07 PS=2.83e-06
mXI58/XI164/XI1/MM0 N_NET069_XI58/XI164/XI1/MM0_d
+ N_XI58/XI164/NET10_XI58/XI164/XI1/MM0_g N_VDD_XI58/XI164/XI1/MM0_s
+ N_VDD_XI32/XI7/MM1_b P_18 L=1.8e-07 W=1.85e-06 AD=4.7175e-13 AS=9.065e-13
+ PD=5.1e-07 PS=2.83e-06
mXI58/XI164/XI1/MM0@2 N_NET069_XI58/XI164/XI1/MM0@2_d
+ N_XI58/XI164/NET10_XI58/XI164/XI1/MM0@2_g N_VDD_XI58/XI164/XI1/MM0@2_s
+ N_VDD_XI32/XI7/MM1_b P_18 L=1.8e-07 W=1.85e-06 AD=4.7175e-13 AS=9.065e-13
+ PD=5.1e-07 PS=2.83e-06
mXI58/XI162/XI0/MM0 N_XI58/XI162/NET8_XI58/XI162/XI0/MM0_d
+ N_NET069_XI58/XI162/XI0/MM0_g N_VDD_XI58/XI162/XI0/MM0_s N_VDD_XI32/XI7/MM1_b
+ P_18 L=1.8e-07 W=1.85e-06 AD=9.065e-13 AS=9.065e-13 PD=2.83e-06 PS=2.83e-06
mXI58/XI162/XI1/MM0 N_XI58/NET086_XI58/XI162/XI1/MM0_d
+ N_XI58/XI162/NET8_XI58/XI162/XI1/MM0_g N_VDD_XI58/XI162/XI1/MM0_s
+ N_VDD_XI32/XI7/MM1_b P_18 L=1.8e-07 W=1.85e-06 AD=9.065e-13 AS=9.065e-13
+ PD=2.83e-06 PS=2.83e-06
mXI58/XI86/XI0/MM0 N_XI58/XI86/NET8_XI58/XI86/XI0/MM0_d
+ N_XI58/NET086_XI58/XI86/XI0/MM0_g N_VDD_XI58/XI86/XI0/MM0_s
+ N_VDD_XI32/XI7/MM1_b P_18 L=1.8e-07 W=1.85e-06 AD=9.065e-13 AS=9.065e-13
+ PD=2.83e-06 PS=2.83e-06
mXI58/XI86/XI1/MM0 N_XI58/NET30_XI58/XI86/XI1/MM0_d
+ N_XI58/XI86/NET8_XI58/XI86/XI1/MM0_g N_VDD_XI58/XI86/XI1/MM0_s
+ N_VDD_XI32/XI7/MM1_b P_18 L=1.8e-07 W=1.85e-06 AD=9.065e-13 AS=9.065e-13
+ PD=2.83e-06 PS=2.83e-06
mXI58/XI99/XI0/MM0 N_XI58/XI99/NET8_XI58/XI99/XI0/MM0_d
+ N_XI58/NET30_XI58/XI99/XI0/MM0_g N_VDD_XI58/XI99/XI0/MM0_s
+ N_VDD_XI32/XI7/MM1_b P_18 L=1.8e-07 W=1.85e-06 AD=9.065e-13 AS=9.065e-13
+ PD=2.83e-06 PS=2.83e-06
mXI58/XI99/XI1/MM0 N_XI58/NET039_XI58/XI99/XI1/MM0_d
+ N_XI58/XI99/NET8_XI58/XI99/XI1/MM0_g N_VDD_XI58/XI99/XI1/MM0_s
+ N_VDD_XI32/XI7/MM1_b P_18 L=1.8e-07 W=1.85e-06 AD=9.065e-13 AS=9.065e-13
+ PD=2.83e-06 PS=2.83e-06
mXI58/XI149/XI0/MM0 N_XI58/XI149/NET8_XI58/XI149/XI0/MM0_d
+ N_XI58/NET039_XI58/XI149/XI0/MM0_g N_VDD_XI58/XI149/XI0/MM0_s
+ N_VDD_XI32/XI7/MM1_b P_18 L=1.8e-07 W=1.85e-06 AD=9.065e-13 AS=9.065e-13
+ PD=2.83e-06 PS=2.83e-06
mXI58/XI149/XI1/MM0 N_XI58/NET081_XI58/XI149/XI1/MM0_d
+ N_XI58/XI149/NET8_XI58/XI149/XI1/MM0_g N_VDD_XI58/XI149/XI1/MM0_s
+ N_VDD_XI32/XI7/MM1_b P_18 L=1.8e-07 W=1.85e-06 AD=9.065e-13 AS=9.065e-13
+ PD=2.83e-06 PS=2.83e-06
mXI58/XI101/XI0/MM0 N_XI58/XI101/NET8_XI58/XI101/XI0/MM0_d
+ N_XI58/NET081_XI58/XI101/XI0/MM0_g N_VDD_XI58/XI101/XI0/MM0_s
+ N_VDD_XI32/XI7/MM1_b P_18 L=1.8e-07 W=1.85e-06 AD=9.065e-13 AS=9.065e-13
+ PD=2.83e-06 PS=2.83e-06
mXI58/XI101/XI1/MM0 N_NET070_XI58/XI101/XI1/MM0_d
+ N_XI58/XI101/NET8_XI58/XI101/XI1/MM0_g N_VDD_XI58/XI101/XI1/MM0_s
+ N_VDD_XI32/XI7/MM1_b P_18 L=1.8e-07 W=1.85e-06 AD=9.065e-13 AS=9.065e-13
+ PD=2.83e-06 PS=2.83e-06
mXI58/XI179/XI0/MM0 N_XI58/XI179/NET10_XI58/XI179/XI0/MM0_d
+ N_NET070_XI58/XI179/XI0/MM0_g N_VDD_XI58/XI179/XI0/MM0_s
+ N_VDD_XI58/XI179/XI0/MM0_b P_18 L=9e-07 W=1.85e-06 AD=2.294e-12 AS=9.065e-13
+ PD=4.33e-06 PS=2.83e-06
mXI58/XI179/XI1/MM0 N_XI58/NET068_XI58/XI179/XI1/MM0_d
+ N_XI58/XI179/NET10_XI58/XI179/XI1/MM0_g N_VDD_XI58/XI179/XI1/MM0_s
+ N_VDD_XI58/XI179/XI0/MM0_b P_18 L=9e-07 W=1.85e-06 AD=2.294e-12 AS=9.065e-13
+ PD=4.33e-06 PS=2.83e-06
mXI58/XI181/XI0/MM0 N_XI58/XI181/NET10_XI58/XI181/XI0/MM0_d
+ N_XI58/NET068_XI58/XI181/XI0/MM0_g N_VDD_XI58/XI181/XI0/MM0_s
+ N_VDD_XI58/XI181/XI0/MM0_b P_18 L=9e-07 W=1.85e-06 AD=2.294e-12 AS=9.065e-13
+ PD=4.33e-06 PS=2.83e-06
mXI58/XI181/XI1/MM0 N_XI58/NET033_XI58/XI181/XI1/MM0_d
+ N_XI58/XI181/NET10_XI58/XI181/XI1/MM0_g N_VDD_XI58/XI181/XI1/MM0_s
+ N_VDD_XI58/XI181/XI0/MM0_b P_18 L=9e-07 W=1.85e-06 AD=2.294e-12 AS=9.065e-13
+ PD=4.33e-06 PS=2.83e-06
mXI58/XI182/XI0/MM0 N_XI58/XI182/NET8_XI58/XI182/XI0/MM0_d
+ N_XI58/NET033_XI58/XI182/XI0/MM0_g N_VDD_XI58/XI182/XI0/MM0_s
+ N_VDD_XI58/XI182/XI0/MM0_b P_18 L=1.8e-07 W=1.85e-06 AD=9.065e-13 AS=9.065e-13
+ PD=2.83e-06 PS=2.83e-06
mXI58/XI182/XI1/MM0 N_XI58/NET049_XI58/XI182/XI1/MM0_d
+ N_XI58/XI182/NET8_XI58/XI182/XI1/MM0_g N_VDD_XI58/XI182/XI1/MM0_s
+ N_VDD_XI58/XI182/XI0/MM0_b P_18 L=1.8e-07 W=1.85e-06 AD=9.065e-13 AS=9.065e-13
+ PD=2.83e-06 PS=2.83e-06
mXI58/XI183/XI0/MM0 N_XI58/XI183/NET8_XI58/XI183/XI0/MM0_d
+ N_XI58/NET049_XI58/XI183/XI0/MM0_g N_VDD_XI58/XI183/XI0/MM0_s
+ N_VDD_XI58/XI182/XI0/MM0_b P_18 L=1.8e-07 W=1.85e-06 AD=9.065e-13 AS=9.065e-13
+ PD=2.83e-06 PS=2.83e-06
mXI58/XI183/XI1/MM0 N_NET068_XI58/XI183/XI1/MM0_d
+ N_XI58/XI183/NET8_XI58/XI183/XI1/MM0_g N_VDD_XI58/XI183/XI1/MM0_s
+ N_VDD_XI58/XI182/XI0/MM0_b P_18 L=1.8e-07 W=1.85e-06 AD=9.065e-13 AS=9.065e-13
+ PD=2.83e-06 PS=2.83e-06
mXI48/XI66/XI5/MM0 N_XI48/XI66/NET21_XI48/XI66/XI5/MM0_d
+ N_XI48/XI66/NET52_XI48/XI66/XI5/MM0_g N_VDD_XI48/XI66/XI5/MM0_s
+ N_VDD_XI48/XI66/MM0_b P_18 L=1.8e-07 W=1.85e-06 AD=9.065e-13 AS=9.065e-13
+ PD=2.83e-06 PS=2.83e-06
mXI48/XI66/XI6/MM0 N_XI48/XI66/NET48_XI48/XI66/XI6/MM0_d
+ N_XI48/XI66/NET21_XI48/XI66/XI6/MM0_g N_VDD_XI48/XI66/XI6/MM0_s
+ N_VDD_XI48/XI66/MM1_b P_18 L=1.8e-07 W=1.85e-06 AD=9.065e-13 AS=9.065e-13
+ PD=2.83e-06 PS=2.83e-06
mXI48/XI65/XI5/MM0 N_XI48/XI65/NET21_XI48/XI65/XI5/MM0_d
+ N_XI48/XI65/NET52_XI48/XI65/XI5/MM0_g N_VDD_XI48/XI65/XI5/MM0_s
+ N_VDD_XI48/XI66/MM1_b P_18 L=1.8e-07 W=1.85e-06 AD=9.065e-13 AS=9.065e-13
+ PD=2.83e-06 PS=2.83e-06
mXI48/XI65/XI6/MM0 N_XI48/XI65/NET48_XI48/XI65/XI6/MM0_d
+ N_XI48/XI65/NET21_XI48/XI65/XI6/MM0_g N_VDD_XI48/XI65/XI6/MM0_s
+ N_VDD_XI48/XI65/MM1_b P_18 L=1.8e-07 W=1.85e-06 AD=9.065e-13 AS=9.065e-13
+ PD=2.83e-06 PS=2.83e-06
mXI48/XI64/XI5/MM0 N_XI48/XI64/NET21_XI48/XI64/XI5/MM0_d
+ N_XI48/XI64/NET52_XI48/XI64/XI5/MM0_g N_VDD_XI48/XI64/XI5/MM0_s
+ N_VDD_XI48/XI65/MM1_b P_18 L=1.8e-07 W=1.85e-06 AD=9.065e-13 AS=9.065e-13
+ PD=2.83e-06 PS=2.83e-06
mXI48/XI64/XI6/MM0 N_XI48/XI64/NET48_XI48/XI64/XI6/MM0_d
+ N_XI48/XI64/NET21_XI48/XI64/XI6/MM0_g N_VDD_XI48/XI64/XI6/MM0_s
+ N_VDD_XI48/XI64/MM1_b P_18 L=1.8e-07 W=1.85e-06 AD=9.065e-13 AS=9.065e-13
+ PD=2.83e-06 PS=2.83e-06
mXI48/XI60/XI6/MM0 N_XI48/XI60/NET48_XI48/XI60/XI6/MM0_d
+ N_XI48/XI60/NET21_XI48/XI60/XI6/MM0_g N_VDD_XI48/XI60/XI6/MM0_s
+ N_VDD_XI48/XI60/MM1_b P_18 L=1.8e-07 W=1.85e-06 AD=9.065e-13 AS=9.065e-13
+ PD=2.83e-06 PS=2.83e-06
mXI48/XI60/XI5/MM0 N_XI48/XI60/NET21_XI48/XI60/XI5/MM0_d
+ N_XI48/XI60/NET52_XI48/XI60/XI5/MM0_g N_VDD_XI48/XI60/XI5/MM0_s
+ N_VDD_XI48/XI60/MM0_b P_18 L=1.8e-07 W=1.85e-06 AD=9.065e-13 AS=9.065e-13
+ PD=2.83e-06 PS=2.83e-06
mXI48/XI61/XI5/MM0 N_XI48/XI61/NET21_XI48/XI61/XI5/MM0_d
+ N_XI48/XI61/NET52_XI48/XI61/XI5/MM0_g N_VDD_XI48/XI61/XI5/MM0_s
+ N_VDD_XI42/XI519/XI72/XI21/MM6_b P_18 L=1.8e-07 W=1.85e-06 AD=9.065e-13
+ AS=9.065e-13 PD=2.83e-06 PS=2.83e-06
mXI48/XI61/XI6/MM0 N_XI48/XI61/NET48_XI48/XI61/XI6/MM0_d
+ N_XI48/XI61/NET21_XI48/XI61/XI6/MM0_g N_VDD_XI48/XI61/XI6/MM0_s
+ N_VDD_XI48/XI61/MM1_b P_18 L=1.8e-07 W=1.85e-06 AD=9.065e-13 AS=9.065e-13
+ PD=2.83e-06 PS=2.83e-06
mXI48/XI62/XI6/MM0 N_XI48/XI62/NET48_XI48/XI62/XI6/MM0_d
+ N_XI48/XI62/NET21_XI48/XI62/XI6/MM0_g N_VDD_XI48/XI62/XI6/MM0_s
+ N_VDD_XI48/XI62/MM1_b P_18 L=1.8e-07 W=1.85e-06 AD=9.065e-13 AS=9.065e-13
+ PD=2.83e-06 PS=2.83e-06
mXI48/XI62/XI5/MM0 N_XI48/XI62/NET21_XI48/XI62/XI5/MM0_d
+ N_XI48/XI62/NET52_XI48/XI62/XI5/MM0_g N_VDD_XI48/XI62/XI5/MM0_s
+ N_VDD_XI48/XI62/MM0_b P_18 L=1.8e-07 W=1.85e-06 AD=9.065e-13 AS=9.065e-13
+ PD=2.83e-06 PS=2.83e-06
mXI48/XI63/XI5/MM0 N_XI48/XI63/NET21_XI48/XI63/XI5/MM0_d
+ N_XI48/XI63/NET52_XI48/XI63/XI5/MM0_g N_VDD_XI48/XI63/XI5/MM0_s
+ N_VDD_XI42/XI519/XI73/XI21/MM6_b P_18 L=1.8e-07 W=1.85e-06 AD=9.065e-13
+ AS=9.065e-13 PD=2.83e-06 PS=2.83e-06
mXI48/XI63/XI6/MM0 N_XI48/XI63/NET48_XI48/XI63/XI6/MM0_d
+ N_XI48/XI63/NET21_XI48/XI63/XI6/MM0_g N_VDD_XI48/XI63/XI6/MM0_s
+ N_VDD_XI48/XI63/MM1_b P_18 L=1.8e-07 W=1.85e-06 AD=9.065e-13 AS=9.065e-13
+ PD=2.83e-06 PS=2.83e-06
mXI32/XI9/XI13/MM0 N_XI32/XI9/NET21_XI32/XI9/XI13/MM0_d
+ N_XI32/XI9/NET52_XI32/XI9/XI13/MM0_g N_VDD_XI32/XI9/XI13/MM0_s
+ N_VDD_XI48/XI63/MM1_b P_18 L=1.8e-07 W=1.85e-06 AD=9.065e-13 AS=9.065e-13
+ PD=2.83e-06 PS=2.83e-06
mXI32/XI9/XI10/MM0 N_XI32/XI9/NET48_XI32/XI9/XI10/MM0_d
+ N_XI32/XI9/NET21_XI32/XI9/XI10/MM0_g N_VDD_XI32/XI9/XI10/MM0_s
+ N_VDD_XI32/XI9/MM1_b P_18 L=1.8e-07 W=1.85e-06 AD=9.065e-13 AS=9.065e-13
+ PD=2.83e-06 PS=2.83e-06
mXI32/XI8/XI13/MM0 N_XI32/XI8/NET21_XI32/XI8/XI13/MM0_d
+ N_XI32/XI8/NET52_XI32/XI8/XI13/MM0_g N_VDD_XI32/XI8/XI13/MM0_s
+ N_VDD_XI32/XI9/MM1_b P_18 L=1.8e-07 W=1.85e-06 AD=9.065e-13 AS=9.065e-13
+ PD=2.83e-06 PS=2.83e-06
mXI32/XI8/XI10/MM0 N_XI32/XI8/NET48_XI32/XI8/XI10/MM0_d
+ N_XI32/XI8/NET21_XI32/XI8/XI10/MM0_g N_VDD_XI32/XI8/XI10/MM0_s
+ N_VDD_XI32/XI8/MM1_b P_18 L=1.8e-07 W=1.85e-06 AD=9.065e-13 AS=9.065e-13
+ PD=2.83e-06 PS=2.83e-06
mXI32/XI7/XI13/MM0 N_XI32/XI7/NET21_XI32/XI7/XI13/MM0_d
+ N_XI32/XI7/NET52_XI32/XI7/XI13/MM0_g N_VDD_XI32/XI7/XI13/MM0_s
+ N_VDD_XI32/XI8/MM1_b P_18 L=1.8e-07 W=1.85e-06 AD=9.065e-13 AS=9.065e-13
+ PD=2.83e-06 PS=2.83e-06
mXI32/XI7/XI10/MM0 N_XI32/XI7/NET48_XI32/XI7/XI10/MM0_d
+ N_XI32/XI7/NET21_XI32/XI7/XI10/MM0_g N_VDD_XI32/XI7/XI10/MM0_s
+ N_VDD_XI32/XI7/MM1_b P_18 L=1.8e-07 W=1.85e-06 AD=9.065e-13 AS=9.065e-13
+ PD=2.83e-06 PS=2.83e-06
mXI42/XI519/XI72/XI20/MM6
+ N_XI42/XI519/XI72/XI20/NET21_XI42/XI519/XI72/XI20/MM6_d
+ N_NET128_XI42/XI519/XI72/XI20/MM6_g N_VDD_XI42/XI519/XI72/XI20/MM6_s
+ N_VDD_XI42/XI519/XI72/XI21/MM6_b P_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13
+ AS=2.632e-13 PD=7.2e-07 PS=1.59e-06
mXI42/XI519/XI73/XI20/MM6
+ N_XI42/XI519/XI73/XI20/NET21_XI42/XI519/XI73/XI20/MM6_d
+ N_NET142_XI42/XI519/XI73/XI20/MM6_g N_VDD_XI42/XI519/XI73/XI20/MM6_s
+ N_VDD_XI42/XI519/XI73/XI21/MM6_b P_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13
+ AS=2.632e-13 PD=7.2e-07 PS=1.59e-06
mXI42/XI519/XI72/XI20/MM7 N_XI42/XI519/NET113_XI42/XI519/XI72/XI20/MM7_d
+ N_NET129_XI42/XI519/XI72/XI20/MM7_g
+ N_XI42/XI519/XI72/XI20/NET21_XI42/XI519/XI72/XI20/MM7_s
+ N_VDD_XI42/XI519/XI72/XI21/MM6_b P_18 L=1.8e-07 W=4.7e-07 AD=2.397e-13
+ AS=1.692e-13 PD=1.49e-06 PS=7.2e-07
mXI42/XI519/XI73/XI20/MM7 N_XI42/XI519/NET31_XI42/XI519/XI73/XI20/MM7_d
+ N_NET143_XI42/XI519/XI73/XI20/MM7_g
+ N_XI42/XI519/XI73/XI20/NET21_XI42/XI519/XI73/XI20/MM7_s
+ N_VDD_XI42/XI519/XI73/XI21/MM6_b P_18 L=1.8e-07 W=4.7e-07 AD=2.397e-13
+ AS=1.692e-13 PD=1.49e-06 PS=7.2e-07
mXI48/XI66/MM2 N_XI48/XI66/NET44_XI48/XI66/MM2_d N_NET90_XI48/XI66/MM2_g
+ N_XI48/XI66/NET21_XI48/XI66/MM2_s N_VDD_XI48/XI66/MM0_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI48/XI66/MM3 N_XI48/XI66/NET059_XI48/XI66/MM3_d N_CLK_XI48/XI66/MM3_g
+ N_XI48/XI66/NET44_XI48/XI66/MM3_s N_VDD_XI48/XI66/MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI48/XI65/MM2 N_XI48/XI65/NET44_XI48/XI65/MM2_d N_NET90_XI48/XI65/MM2_g
+ N_XI48/XI65/NET21_XI48/XI65/MM2_s N_VDD_XI48/XI66/MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI48/XI65/MM3 N_XI48/XI65/NET059_XI48/XI65/MM3_d N_CLK_XI48/XI65/MM3_g
+ N_XI48/XI65/NET44_XI48/XI65/MM3_s N_VDD_XI48/XI65/MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI48/XI64/MM2 N_XI48/XI64/NET44_XI48/XI64/MM2_d N_NET90_XI48/XI64/MM2_g
+ N_XI48/XI64/NET21_XI48/XI64/MM2_s N_VDD_XI48/XI65/MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI48/XI64/MM3 N_XI48/XI64/NET059_XI48/XI64/MM3_d N_CLK_XI48/XI64/MM3_g
+ N_XI48/XI64/NET44_XI48/XI64/MM3_s N_VDD_XI48/XI64/MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI48/XI60/MM3 N_XI48/XI60/NET059_XI48/XI60/MM3_d N_CLK_XI48/XI60/MM3_g
+ N_XI48/XI60/NET44_XI48/XI60/MM3_s N_VDD_XI48/XI60/MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI48/XI60/MM2 N_XI48/XI60/NET44_XI48/XI60/MM2_d N_NET90_XI48/XI60/MM2_g
+ N_XI48/XI60/NET21_XI48/XI60/MM2_s N_VDD_XI48/XI60/MM0_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI48/XI61/MM2 N_XI48/XI61/NET44_XI48/XI61/MM2_d N_NET90_XI48/XI61/MM2_g
+ N_XI48/XI61/NET21_XI48/XI61/MM2_s N_VDD_XI42/XI519/XI72/XI21/MM6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI48/XI61/MM3 N_XI48/XI61/NET059_XI48/XI61/MM3_d N_CLK_XI48/XI61/MM3_g
+ N_XI48/XI61/NET44_XI48/XI61/MM3_s N_VDD_XI48/XI61/MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI48/XI62/MM3 N_XI48/XI62/NET059_XI48/XI62/MM3_d N_CLK_XI48/XI62/MM3_g
+ N_XI48/XI62/NET44_XI48/XI62/MM3_s N_VDD_XI48/XI62/MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI48/XI62/MM2 N_XI48/XI62/NET44_XI48/XI62/MM2_d N_NET90_XI48/XI62/MM2_g
+ N_XI48/XI62/NET21_XI48/XI62/MM2_s N_VDD_XI48/XI62/MM0_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI48/XI63/MM2 N_XI48/XI63/NET44_XI48/XI63/MM2_d N_NET90_XI48/XI63/MM2_g
+ N_XI48/XI63/NET21_XI48/XI63/MM2_s N_VDD_XI42/XI519/XI73/XI21/MM6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI48/XI63/MM3 N_XI48/XI63/NET059_XI48/XI63/MM3_d N_CLK_XI48/XI63/MM3_g
+ N_XI48/XI63/NET44_XI48/XI63/MM3_s N_VDD_XI48/XI63/MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI32/XI9/MM2 N_XI32/XI9/NET44_XI32/XI9/MM2_d N_NET90_XI32/XI9/MM2_g
+ N_XI32/XI9/NET21_XI32/XI9/MM2_s N_VDD_XI48/XI63/MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI32/XI9/MM3 N_NET434_XI32/XI9/MM3_d N_CLK_XI32/XI9/MM3_g
+ N_XI32/XI9/NET44_XI32/XI9/MM3_s N_VDD_XI32/XI9/MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI32/XI8/MM2 N_XI32/XI8/NET44_XI32/XI8/MM2_d N_NET90_XI32/XI8/MM2_g
+ N_XI32/XI8/NET21_XI32/XI8/MM2_s N_VDD_XI32/XI9/MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI32/XI8/MM3 N_NET435_XI32/XI8/MM3_d N_CLK_XI32/XI8/MM3_g
+ N_XI32/XI8/NET44_XI32/XI8/MM3_s N_VDD_XI32/XI8/MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI32/XI7/MM2 N_XI32/XI7/NET44_XI32/XI7/MM2_d N_NET90_XI32/XI7/MM2_g
+ N_XI32/XI7/NET21_XI32/XI7/MM2_s N_VDD_XI32/XI8/MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI32/XI7/MM3 N_NET436_XI32/XI7/MM3_d N_CLK_XI32/XI7/MM3_g
+ N_XI32/XI7/NET44_XI32/XI7/MM3_s N_VDD_XI32/XI7/MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI42/XI519/XI72/XI19/MM6
+ N_XI42/XI519/XI72/XI19/NET21_XI42/XI519/XI72/XI19/MM6_d
+ N_NET127_XI42/XI519/XI72/XI19/MM6_g N_VDD_XI42/XI519/XI72/XI19/MM6_s
+ N_VDD_XI42/XI519/XI72/XI21/MM6_b P_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13
+ AS=2.632e-13 PD=7.2e-07 PS=1.59e-06
mXI42/XI519/XI73/XI19/MM6
+ N_XI42/XI519/XI73/XI19/NET21_XI42/XI519/XI73/XI19/MM6_d
+ N_NET141_XI42/XI519/XI73/XI19/MM6_g N_VDD_XI42/XI519/XI73/XI19/MM6_s
+ N_VDD_XI42/XI519/XI73/XI21/MM6_b P_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13
+ AS=2.632e-13 PD=7.2e-07 PS=1.59e-06
mXI48/XI66/XI7/MM0 N_XI48/NET0110_XI48/XI66/XI7/MM0_d
+ N_XI48/XI66/NET44_XI48/XI66/XI7/MM0_g N_VDD_XI48/XI66/XI7/MM0_s
+ N_VDD_XI48/XI66/MM0_b P_18 L=1.8e-07 W=1.85e-06 AD=9.065e-13 AS=9.065e-13
+ PD=2.83e-06 PS=2.83e-06
mXI48/XI66/XI8/MM0 N_XI48/XI66/NET059_XI48/XI66/XI8/MM0_d
+ N_XI48/NET0110_XI48/XI66/XI8/MM0_g N_VDD_XI48/XI66/XI8/MM0_s
+ N_VDD_XI48/XI66/MM1_b P_18 L=1.8e-07 W=1.85e-06 AD=9.065e-13 AS=9.065e-13
+ PD=2.83e-06 PS=2.83e-06
mXI48/XI65/XI7/MM0 N_XI48/NET098_XI48/XI65/XI7/MM0_d
+ N_XI48/XI65/NET44_XI48/XI65/XI7/MM0_g N_VDD_XI48/XI65/XI7/MM0_s
+ N_VDD_XI48/XI66/MM1_b P_18 L=1.8e-07 W=1.85e-06 AD=9.065e-13 AS=9.065e-13
+ PD=2.83e-06 PS=2.83e-06
mXI48/XI65/XI8/MM0 N_XI48/XI65/NET059_XI48/XI65/XI8/MM0_d
+ N_XI48/NET098_XI48/XI65/XI8/MM0_g N_VDD_XI48/XI65/XI8/MM0_s
+ N_VDD_XI48/XI65/MM1_b P_18 L=1.8e-07 W=1.85e-06 AD=9.065e-13 AS=9.065e-13
+ PD=2.83e-06 PS=2.83e-06
mXI48/XI64/XI7/MM0 N_XI48/NET0116_XI48/XI64/XI7/MM0_d
+ N_XI48/XI64/NET44_XI48/XI64/XI7/MM0_g N_VDD_XI48/XI64/XI7/MM0_s
+ N_VDD_XI48/XI65/MM1_b P_18 L=1.8e-07 W=1.85e-06 AD=9.065e-13 AS=9.065e-13
+ PD=2.83e-06 PS=2.83e-06
mXI48/XI64/XI8/MM0 N_XI48/XI64/NET059_XI48/XI64/XI8/MM0_d
+ N_XI48/NET0116_XI48/XI64/XI8/MM0_g N_VDD_XI48/XI64/XI8/MM0_s
+ N_VDD_XI48/XI64/MM1_b P_18 L=1.8e-07 W=1.85e-06 AD=9.065e-13 AS=9.065e-13
+ PD=2.83e-06 PS=2.83e-06
mXI48/XI60/XI8/MM0 N_XI48/XI60/NET059_XI48/XI60/XI8/MM0_d
+ N_XI48/NET0122_XI48/XI60/XI8/MM0_g N_VDD_XI48/XI60/XI8/MM0_s
+ N_VDD_XI48/XI60/MM1_b P_18 L=1.8e-07 W=1.85e-06 AD=9.065e-13 AS=9.065e-13
+ PD=2.83e-06 PS=2.83e-06
mXI48/XI60/XI7/MM0 N_XI48/NET0122_XI48/XI60/XI7/MM0_d
+ N_XI48/XI60/NET44_XI48/XI60/XI7/MM0_g N_VDD_XI48/XI60/XI7/MM0_s
+ N_VDD_XI48/XI60/MM0_b P_18 L=1.8e-07 W=1.85e-06 AD=9.065e-13 AS=9.065e-13
+ PD=2.83e-06 PS=2.83e-06
mXI48/XI61/XI7/MM0 N_XI48/NET0134_XI48/XI61/XI7/MM0_d
+ N_XI48/XI61/NET44_XI48/XI61/XI7/MM0_g N_VDD_XI48/XI61/XI7/MM0_s
+ N_VDD_XI42/XI519/XI72/XI21/MM6_b P_18 L=1.8e-07 W=1.85e-06 AD=9.065e-13
+ AS=9.065e-13 PD=2.83e-06 PS=2.83e-06
mXI48/XI61/XI8/MM0 N_XI48/XI61/NET059_XI48/XI61/XI8/MM0_d
+ N_XI48/NET0134_XI48/XI61/XI8/MM0_g N_VDD_XI48/XI61/XI8/MM0_s
+ N_VDD_XI48/XI61/MM1_b P_18 L=1.8e-07 W=1.85e-06 AD=9.065e-13 AS=9.065e-13
+ PD=2.83e-06 PS=2.83e-06
mXI48/XI62/XI8/MM0 N_XI48/XI62/NET059_XI48/XI62/XI8/MM0_d
+ N_XI48/NET0128_XI48/XI62/XI8/MM0_g N_VDD_XI48/XI62/XI8/MM0_s
+ N_VDD_XI48/XI62/MM1_b P_18 L=1.8e-07 W=1.85e-06 AD=9.065e-13 AS=9.065e-13
+ PD=2.83e-06 PS=2.83e-06
mXI48/XI62/XI7/MM0 N_XI48/NET0128_XI48/XI62/XI7/MM0_d
+ N_XI48/XI62/NET44_XI48/XI62/XI7/MM0_g N_VDD_XI48/XI62/XI7/MM0_s
+ N_VDD_XI48/XI62/MM0_b P_18 L=1.8e-07 W=1.85e-06 AD=9.065e-13 AS=9.065e-13
+ PD=2.83e-06 PS=2.83e-06
mXI48/XI63/XI7/MM0 N_XI48/NET0104_XI48/XI63/XI7/MM0_d
+ N_XI48/XI63/NET44_XI48/XI63/XI7/MM0_g N_VDD_XI48/XI63/XI7/MM0_s
+ N_VDD_XI42/XI519/XI73/XI21/MM6_b P_18 L=1.8e-07 W=1.85e-06 AD=9.065e-13
+ AS=9.065e-13 PD=2.83e-06 PS=2.83e-06
mXI48/XI63/XI8/MM0 N_XI48/XI63/NET059_XI48/XI63/XI8/MM0_d
+ N_XI48/NET0104_XI48/XI63/XI8/MM0_g N_VDD_XI48/XI63/XI8/MM0_s
+ N_VDD_XI48/XI63/MM1_b P_18 L=1.8e-07 W=1.85e-06 AD=9.065e-13 AS=9.065e-13
+ PD=2.83e-06 PS=2.83e-06
mXI32/XI9/XI12/MM0 N_NET437_XI32/XI9/XI12/MM0_d
+ N_XI32/XI9/NET44_XI32/XI9/XI12/MM0_g N_VDD_XI32/XI9/XI12/MM0_s
+ N_VDD_XI48/XI63/MM1_b P_18 L=1.8e-07 W=1.85e-06 AD=9.065e-13 AS=9.065e-13
+ PD=2.83e-06 PS=2.83e-06
mXI32/XI9/XI11/MM0 N_NET434_XI32/XI9/XI11/MM0_d N_NET437_XI32/XI9/XI11/MM0_g
+ N_VDD_XI32/XI9/XI11/MM0_s N_VDD_XI32/XI9/MM1_b P_18 L=1.8e-07 W=1.85e-06
+ AD=9.065e-13 AS=9.065e-13 PD=2.83e-06 PS=2.83e-06
mXI32/XI8/XI12/MM0 N_NET438_XI32/XI8/XI12/MM0_d
+ N_XI32/XI8/NET44_XI32/XI8/XI12/MM0_g N_VDD_XI32/XI8/XI12/MM0_s
+ N_VDD_XI32/XI9/MM1_b P_18 L=1.8e-07 W=1.85e-06 AD=9.065e-13 AS=9.065e-13
+ PD=2.83e-06 PS=2.83e-06
mXI32/XI8/XI11/MM0 N_NET435_XI32/XI8/XI11/MM0_d N_NET438_XI32/XI8/XI11/MM0_g
+ N_VDD_XI32/XI8/XI11/MM0_s N_VDD_XI32/XI8/MM1_b P_18 L=1.8e-07 W=1.85e-06
+ AD=9.065e-13 AS=9.065e-13 PD=2.83e-06 PS=2.83e-06
mXI32/XI7/XI12/MM0 N_NET439_XI32/XI7/XI12/MM0_d
+ N_XI32/XI7/NET44_XI32/XI7/XI12/MM0_g N_VDD_XI32/XI7/XI12/MM0_s
+ N_VDD_XI32/XI8/MM1_b P_18 L=1.8e-07 W=1.85e-06 AD=9.065e-13 AS=9.065e-13
+ PD=2.83e-06 PS=2.83e-06
mXI32/XI7/XI11/MM0 N_NET436_XI32/XI7/XI11/MM0_d N_NET439_XI32/XI7/XI11/MM0_g
+ N_VDD_XI32/XI7/XI11/MM0_s N_VDD_XI32/XI7/MM1_b P_18 L=1.8e-07 W=1.85e-06
+ AD=9.065e-13 AS=9.065e-13 PD=2.83e-06 PS=2.83e-06
mXI42/XI519/XI72/XI19/MM7 N_XI42/XI519/NET112_XI42/XI519/XI72/XI19/MM7_d
+ N_NET130_XI42/XI519/XI72/XI19/MM7_g
+ N_XI42/XI519/XI72/XI19/NET21_XI42/XI519/XI72/XI19/MM7_s
+ N_VDD_XI42/XI519/XI72/XI21/MM6_b P_18 L=1.8e-07 W=4.7e-07 AD=2.397e-13
+ AS=1.692e-13 PD=1.49e-06 PS=7.2e-07
mXI42/XI519/XI73/XI19/MM7 N_XI42/XI519/NET104_XI42/XI519/XI73/XI19/MM7_d
+ N_NET126_XI42/XI519/XI73/XI19/MM7_g
+ N_XI42/XI519/XI73/XI19/NET21_XI42/XI519/XI73/XI19/MM7_s
+ N_VDD_XI42/XI519/XI73/XI21/MM6_b P_18 L=1.8e-07 W=4.7e-07 AD=2.397e-13
+ AS=1.692e-13 PD=1.49e-06 PS=7.2e-07
mXI48/XI68/XI3/MM0 N_NET130_XI48/XI68/XI3/MM0_d N_NET129_XI48/XI68/XI3/MM0_g
+ N_VDD_XI48/XI68/XI3/MM0_s N_VDD_XI48/XI60/MM0_b P_18 L=1.8e-07 W=1.85e-06
+ AD=9.435e-13 AS=9.435e-13 PD=2.87e-06 PS=2.87e-06
mXI48/XI69/XI3/MM0 N_NET128_XI48/XI69/XI3/MM0_d N_NET127_XI48/XI69/XI3/MM0_g
+ N_VDD_XI48/XI69/XI3/MM0_s N_VDD_XI42/XI519/XI72/XI21/MM6_b P_18 L=1.8e-07
+ W=1.85e-06 AD=9.435e-13 AS=9.435e-13 PD=2.87e-06 PS=2.87e-06
mXI48/XI70/XI3/MM0 N_NET126_XI48/XI70/XI3/MM0_d N_NET143_XI48/XI70/XI3/MM0_g
+ N_VDD_XI48/XI70/XI3/MM0_s N_VDD_XI48/XI62/MM0_b P_18 L=1.8e-07 W=1.85e-06
+ AD=9.435e-13 AS=9.435e-13 PD=2.87e-06 PS=2.87e-06
mXI48/XI71/XI3/MM0 N_NET142_XI48/XI71/XI3/MM0_d N_NET141_XI48/XI71/XI3/MM0_g
+ N_VDD_XI48/XI71/XI3/MM0_s N_VDD_XI42/XI519/XI73/XI21/MM6_b P_18 L=1.8e-07
+ W=1.85e-06 AD=9.435e-13 AS=9.435e-13 PD=2.87e-06 PS=2.87e-06
mXI42/XI652/XI0/MM0 N_XI42/XI652/NET8_XI42/XI652/XI0/MM0_d
+ N_XI42/NET01023_XI42/XI652/XI0/MM0_g N_VDD_XI42/XI652/XI0/MM0_s
+ N_VDD_XI48/XI66/MM0_b P_18 L=1.8e-07 W=1.85e-06 AD=9.065e-13 AS=9.065e-13
+ PD=2.83e-06 PS=2.83e-06
mXI48/XI74/XI2/MM1 N_NET135_XI48/XI74/XI2/MM1_d
+ N_XI48/NET0110_XI48/XI74/XI2/MM1_g N_VDD_XI48/XI74/XI2/MM1_s
+ N_VDD_XI48/XI66/MM1_b P_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13 AS=2.632e-13
+ PD=7.2e-07 PS=1.59e-06
mXI48/XI73/XI2/MM1 N_NET137_XI48/XI73/XI2/MM1_d
+ N_XI48/NET098_XI48/XI73/XI2/MM1_g N_VDD_XI48/XI73/XI2/MM1_s
+ N_VDD_XI48/XI66/MM1_b P_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13 AS=2.632e-13
+ PD=7.2e-07 PS=1.59e-06
mXI48/XI72/XI2/MM1 N_NET139_XI48/XI72/XI2/MM1_d
+ N_XI48/NET0116_XI48/XI72/XI2/MM1_g N_VDD_XI48/XI72/XI2/MM1_s
+ N_VDD_XI48/XI65/MM1_b P_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13 AS=2.632e-13
+ PD=7.2e-07 PS=1.59e-06
mXI42/XI519/XI72/XI18/MM6
+ N_XI42/XI519/XI72/XI18/NET21_XI42/XI519/XI72/XI18/MM6_d
+ N_NET128_XI42/XI519/XI72/XI18/MM6_g N_VDD_XI42/XI519/XI72/XI18/MM6_s
+ N_VDD_XI42/XI519/XI72/XI21/MM6_b P_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13
+ AS=2.632e-13 PD=7.2e-07 PS=1.59e-06
mXI42/XI519/XI73/XI18/MM6
+ N_XI42/XI519/XI73/XI18/NET21_XI42/XI519/XI73/XI18/MM6_d
+ N_NET142_XI42/XI519/XI73/XI18/MM6_g N_VDD_XI42/XI519/XI73/XI18/MM6_s
+ N_VDD_XI42/XI519/XI73/XI21/MM6_b P_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13
+ AS=2.632e-13 PD=7.2e-07 PS=1.59e-06
mXI48/XI69/XI2/MM0 N_NET127_XI48/XI69/XI2/MM0_d N_NET069_XI48/XI69/XI2/MM0_g
+ N_VDD_XI48/XI69/XI2/MM0_s N_VDD_XI42/XI519/XI72/XI21/MM6_b P_18 L=1.8e-07
+ W=4.7e-07 AD=1.692e-13 AS=2.397e-13 PD=7.2e-07 PS=1.49e-06
mXI48/XI69/XI2/MM1 N_NET127_XI48/XI69/XI2/MM1_d
+ N_XI48/NET0134_XI48/XI69/XI2/MM1_g N_VDD_XI48/XI69/XI2/MM1_s
+ N_VDD_XI42/XI519/XI72/XI21/MM6_b P_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13
+ AS=2.632e-13 PD=7.2e-07 PS=1.59e-06
mXI48/XI71/XI2/MM0 N_NET141_XI48/XI71/XI2/MM0_d N_NET069_XI48/XI71/XI2/MM0_g
+ N_VDD_XI48/XI71/XI2/MM0_s N_VDD_XI42/XI519/XI73/XI21/MM6_b P_18 L=1.8e-07
+ W=4.7e-07 AD=1.692e-13 AS=2.397e-13 PD=7.2e-07 PS=1.49e-06
mXI48/XI71/XI2/MM1 N_NET141_XI48/XI71/XI2/MM1_d
+ N_XI48/NET0104_XI48/XI71/XI2/MM1_g N_VDD_XI48/XI71/XI2/MM1_s
+ N_VDD_XI42/XI519/XI73/XI21/MM6_b P_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13
+ AS=2.632e-13 PD=7.2e-07 PS=1.59e-06
mXI48/XI68/XI2/MM1 N_NET129_XI48/XI68/XI2/MM1_d
+ N_XI48/NET0122_XI48/XI68/XI2/MM1_g N_VDD_XI48/XI68/XI2/MM1_s
+ N_VDD_XI48/XI60/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13 AS=2.632e-13
+ PD=7.2e-07 PS=1.59e-06
mXI48/XI68/XI2/MM0 N_NET129_XI48/XI68/XI2/MM0_d N_NET069_XI48/XI68/XI2/MM0_g
+ N_VDD_XI48/XI68/XI2/MM0_s N_VDD_XI48/XI60/MM0_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.692e-13 AS=2.397e-13 PD=7.2e-07 PS=1.49e-06
mXI48/XI70/XI2/MM1 N_NET143_XI48/XI70/XI2/MM1_d
+ N_XI48/NET0128_XI48/XI70/XI2/MM1_g N_VDD_XI48/XI70/XI2/MM1_s
+ N_VDD_XI48/XI62/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13 AS=2.632e-13
+ PD=7.2e-07 PS=1.59e-06
mXI48/XI70/XI2/MM0 N_NET143_XI48/XI70/XI2/MM0_d N_NET069_XI48/XI70/XI2/MM0_g
+ N_VDD_XI48/XI70/XI2/MM0_s N_VDD_XI48/XI62/MM0_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.692e-13 AS=2.397e-13 PD=7.2e-07 PS=1.49e-06
mXI48/XI74/XI2/MM0 N_NET135_XI48/XI74/XI2/MM0_d N_NET069_XI48/XI74/XI2/MM0_g
+ N_VDD_XI48/XI74/XI2/MM0_s N_VDD_XI48/XI66/MM1_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.692e-13 AS=2.397e-13 PD=7.2e-07 PS=1.49e-06
mXI48/XI73/XI2/MM0 N_NET137_XI48/XI73/XI2/MM0_d N_NET069_XI48/XI73/XI2/MM0_g
+ N_VDD_XI48/XI73/XI2/MM0_s N_VDD_XI48/XI66/MM1_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.692e-13 AS=2.397e-13 PD=7.2e-07 PS=1.49e-06
mXI48/XI72/XI2/MM0 N_NET139_XI48/XI72/XI2/MM0_d N_NET069_XI48/XI72/XI2/MM0_g
+ N_VDD_XI48/XI72/XI2/MM0_s N_VDD_XI48/XI65/MM1_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.692e-13 AS=2.397e-13 PD=7.2e-07 PS=1.49e-06
mXI42/XI519/XI72/XI18/MM7 N_XI42/XI519/NET111_XI42/XI519/XI72/XI18/MM7_d
+ N_NET130_XI42/XI519/XI72/XI18/MM7_g
+ N_XI42/XI519/XI72/XI18/NET21_XI42/XI519/XI72/XI18/MM7_s
+ N_VDD_XI42/XI519/XI72/XI21/MM6_b P_18 L=1.8e-07 W=4.7e-07 AD=2.397e-13
+ AS=1.692e-13 PD=1.49e-06 PS=7.2e-07
mXI42/XI519/XI73/XI18/MM7 N_XI42/XI519/NET103_XI42/XI519/XI73/XI18/MM7_d
+ N_NET126_XI42/XI519/XI73/XI18/MM7_g
+ N_XI42/XI519/XI73/XI18/NET21_XI42/XI519/XI73/XI18/MM7_s
+ N_VDD_XI42/XI519/XI73/XI21/MM6_b P_18 L=1.8e-07 W=4.7e-07 AD=2.397e-13
+ AS=1.692e-13 PD=1.49e-06 PS=7.2e-07
mXI30/XI67/MM2 N_NET470_XI30/XI67/MM2_d N_NET437_XI30/XI67/MM2_g
+ N_VDD_XI30/XI67/MM2_s N_VDD_XI30/XI67/MM2_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI30/XI67/MM1 N_NET470_XI30/XI67/MM1_d N_NET438_XI30/XI67/MM1_g
+ N_VDD_XI30/XI67/MM1_s N_VDD_XI30/XI67/MM2_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI30/XI67/MM0 N_NET470_XI30/XI67/MM0_d N_NET439_XI30/XI67/MM0_g
+ N_VDD_XI30/XI67/MM0_s N_VDD_XI30/XI67/MM2_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI30/XI69/MM2 N_NET468_XI30/XI69/MM2_d N_NET437_XI30/XI69/MM2_g
+ N_VDD_XI30/XI69/MM2_s N_VDD_XI30/XI67/MM2_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI30/XI69/MM1 N_NET468_XI30/XI69/MM1_d N_NET435_XI30/XI69/MM1_g
+ N_VDD_XI30/XI69/MM1_s N_VDD_XI30/XI67/MM2_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI30/XI69/MM0 N_NET468_XI30/XI69/MM0_d N_NET439_XI30/XI69/MM0_g
+ N_VDD_XI30/XI69/MM0_s N_VDD_XI30/XI67/MM2_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI30/XI71/MM2 N_NET466_XI30/XI71/MM2_d N_NET437_XI30/XI71/MM2_g
+ N_VDD_XI30/XI71/MM2_s N_VDD_XI30/XI67/MM2_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI30/XI71/MM1 N_NET466_XI30/XI71/MM1_d N_NET438_XI30/XI71/MM1_g
+ N_VDD_XI30/XI71/MM1_s N_VDD_XI30/XI67/MM2_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI30/XI71/MM0 N_NET466_XI30/XI71/MM0_d N_NET436_XI30/XI71/MM0_g
+ N_VDD_XI30/XI71/MM0_s N_VDD_XI30/XI67/MM2_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI30/XI73/MM2 N_NET464_XI30/XI73/MM2_d N_NET437_XI30/XI73/MM2_g
+ N_VDD_XI30/XI73/MM2_s N_VDD_XI30/XI67/MM2_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI30/XI73/MM1 N_NET464_XI30/XI73/MM1_d N_NET435_XI30/XI73/MM1_g
+ N_VDD_XI30/XI73/MM1_s N_VDD_XI30/XI67/MM2_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI30/XI73/MM0 N_NET464_XI30/XI73/MM0_d N_NET436_XI30/XI73/MM0_g
+ N_VDD_XI30/XI73/MM0_s N_VDD_XI30/XI67/MM2_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI30/XI68/MM2 N_NET469_XI30/XI68/MM2_d N_NET434_XI30/XI68/MM2_g
+ N_VDD_XI30/XI68/MM2_s N_VDD_XI30/XI67/MM2_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI30/XI68/MM1 N_NET469_XI30/XI68/MM1_d N_NET438_XI30/XI68/MM1_g
+ N_VDD_XI30/XI68/MM1_s N_VDD_XI30/XI67/MM2_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI30/XI68/MM0 N_NET469_XI30/XI68/MM0_d N_NET439_XI30/XI68/MM0_g
+ N_VDD_XI30/XI68/MM0_s N_VDD_XI30/XI67/MM2_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI30/XI70/MM2 N_NET467_XI30/XI70/MM2_d N_NET434_XI30/XI70/MM2_g
+ N_VDD_XI30/XI70/MM2_s N_VDD_XI30/XI67/MM2_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI30/XI70/MM1 N_NET467_XI30/XI70/MM1_d N_NET435_XI30/XI70/MM1_g
+ N_VDD_XI30/XI70/MM1_s N_VDD_XI30/XI67/MM2_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI30/XI70/MM0 N_NET467_XI30/XI70/MM0_d N_NET439_XI30/XI70/MM0_g
+ N_VDD_XI30/XI70/MM0_s N_VDD_XI30/XI67/MM2_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI30/XI72/MM2 N_NET465_XI30/XI72/MM2_d N_NET434_XI30/XI72/MM2_g
+ N_VDD_XI30/XI72/MM2_s N_VDD_XI30/XI67/MM2_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI30/XI72/MM1 N_NET465_XI30/XI72/MM1_d N_NET438_XI30/XI72/MM1_g
+ N_VDD_XI30/XI72/MM1_s N_VDD_XI30/XI67/MM2_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI30/XI72/MM0 N_NET465_XI30/XI72/MM0_d N_NET436_XI30/XI72/MM0_g
+ N_VDD_XI30/XI72/MM0_s N_VDD_XI30/XI67/MM2_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI30/XI74/MM2 N_NET463_XI30/XI74/MM2_d N_NET434_XI30/XI74/MM2_g
+ N_VDD_XI30/XI74/MM2_s N_VDD_XI30/XI67/MM2_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI30/XI74/MM1 N_NET463_XI30/XI74/MM1_d N_NET435_XI30/XI74/MM1_g
+ N_VDD_XI30/XI74/MM1_s N_VDD_XI30/XI67/MM2_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI30/XI74/MM0 N_NET463_XI30/XI74/MM0_d N_NET436_XI30/XI74/MM0_g
+ N_VDD_XI30/XI74/MM0_s N_VDD_XI30/XI67/MM2_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI42/XI652/XI1/MM0 N_NET0133_XI42/XI652/XI1/MM0_d
+ N_XI42/XI652/NET8_XI42/XI652/XI1/MM0_g N_VDD_XI42/XI652/XI1/MM0_s
+ N_VDD_XI48/XI66/MM0_b P_18 L=1.8e-07 W=1.85e-06 AD=9.065e-13 AS=9.065e-13
+ PD=2.83e-06 PS=2.83e-06
mXI54/XI0/XI10/MM7 N_DOUT<0>_XI54/XI0/XI10/MM7_d
+ N_XI54/NET10_XI54/XI0/XI10/MM7_g N_XI54/XI0/XI10/NET21_XI54/XI0/XI10/MM7_s
+ N_VDD_XI30/XI67/MM2_b P_18 L=1.8e-07 W=4.7e-07 AD=2.3265e-13 AS=1.68025e-13
+ PD=1.46e-06 PS=7.15e-07
mXI54/XI0/XI9/MM7 N_XI54/NET10_XI54/XI0/XI9/MM7_d
+ N_XI54/XI0/NET10_XI54/XI0/XI9/MM7_g N_XI54/XI0/XI9/NET21_XI54/XI0/XI9/MM7_s
+ N_VDD_XI30/XI67/MM2_b P_18 L=1.8e-07 W=4.7e-07 AD=2.3265e-13 AS=1.68025e-13
+ PD=1.46e-06 PS=7.15e-07
mXI54/XI0/XI10/MM6 N_XI54/XI0/XI10/NET21_XI54/XI0/XI10/MM6_d
+ N_XI54/XI0/NET9_XI54/XI0/XI10/MM6_g N_VDD_XI54/XI0/XI10/MM6_s
+ N_VDD_XI30/XI67/MM2_b P_18 L=1.8e-07 W=4.7e-07 AD=1.68025e-13 AS=2.303e-13
+ PD=7.15e-07 PS=1.45e-06
mXI54/XI0/XI9/MM6 N_XI54/XI0/XI9/NET21_XI54/XI0/XI9/MM6_d
+ N_DOUT<0>_XI54/XI0/XI9/MM6_g N_VDD_XI54/XI0/XI9/MM6_s N_VDD_XI30/XI67/MM2_b
+ P_18 L=1.8e-07 W=4.7e-07 AD=1.68025e-13 AS=2.5145e-13 PD=7.15e-07 PS=1.54e-06
mXI54/XI0/XI8/XI2/MM0 N_XI54/XI0/NET9_XI54/XI0/XI8/XI2/MM0_d
+ N_XI54/XI0/XI8/NET12_XI54/XI0/XI8/XI2/MM0_g N_VDD_XI54/XI0/XI8/XI2/MM0_s
+ N_VDD_XI30/XI67/MM2_b P_18 L=1.8e-07 W=1.85e-06 AD=9.435e-13 AS=9.435e-13
+ PD=2.87e-06 PS=2.87e-06
mXI54/XI0/XI7/XI2/MM0 N_XI54/XI0/NET10_XI54/XI0/XI7/XI2/MM0_d
+ N_XI54/XI0/XI7/NET12_XI54/XI0/XI7/XI2/MM0_g N_VDD_XI54/XI0/XI7/XI2/MM0_s
+ N_VDD_XI30/XI67/MM2_b P_18 L=1.8e-07 W=1.85e-06 AD=9.435e-13 AS=9.435e-13
+ PD=2.87e-06 PS=2.87e-06
mXI54/XI0/XI8/XI3/MM0 N_XI54/XI0/XI8/NET12_XI54/XI0/XI8/XI3/MM0_d
+ N_NET068_XI54/XI0/XI8/XI3/MM0_g N_VDD_XI54/XI0/XI8/XI3/MM0_s
+ N_VDD_XI30/XI67/MM2_b P_18 L=1.8e-07 W=4.7e-07 AD=1.68025e-13 AS=2.3265e-13
+ PD=7.15e-07 PS=1.46e-06
mXI54/XI0/XI7/XI3/MM0 N_XI54/XI0/XI7/NET12_XI54/XI0/XI7/XI3/MM0_d
+ N_NET068_XI54/XI0/XI7/XI3/MM0_g N_VDD_XI54/XI0/XI7/XI3/MM0_s
+ N_VDD_XI30/XI67/MM2_b P_18 L=1.8e-07 W=4.7e-07 AD=1.68025e-13 AS=2.3265e-13
+ PD=7.15e-07 PS=1.46e-06
mXI42/XI519/XI86/MM0 N_XI42/NET780_XI42/XI519/XI86/MM0_d
+ N_XI42/XI519/NET114_XI42/XI519/XI86/MM0_g N_VDD_XI42/XI519/XI86/MM0_s
+ N_VDD_XI42/XI519/XI86/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13 AS=2.397e-13
+ PD=7.2e-07 PS=1.49e-06
mXI42/XI519/XI86/MM1 N_XI42/NET780_XI42/XI519/XI86/MM1_d
+ N_XI42/XI519/NET36_XI42/XI519/XI86/MM1_g N_VDD_XI42/XI519/XI86/MM1_s
+ N_VDD_XI42/XI519/XI86/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13 AS=2.632e-13
+ PD=7.2e-07 PS=1.59e-06
mXI42/XI519/XI87/MM0 N_XI42/NET781_XI42/XI519/XI87/MM0_d
+ N_XI42/XI519/NET114_XI42/XI519/XI87/MM0_g N_VDD_XI42/XI519/XI87/MM0_s
+ N_VDD_XI42/XI519/XI87/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13 AS=2.397e-13
+ PD=7.2e-07 PS=1.49e-06
mXI42/XI519/XI87/MM1 N_XI42/NET781_XI42/XI519/XI87/MM1_d
+ N_XI42/XI519/NET31_XI42/XI519/XI87/MM1_g N_VDD_XI42/XI519/XI87/MM1_s
+ N_VDD_XI42/XI519/XI87/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13 AS=2.632e-13
+ PD=7.2e-07 PS=1.59e-06
mXI42/XI519/XI88/MM0 N_XI42/NET782_XI42/XI519/XI88/MM0_d
+ N_XI42/XI519/NET114_XI42/XI519/XI88/MM0_g N_VDD_XI42/XI519/XI88/MM0_s
+ N_VDD_XI42/XI519/XI88/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13 AS=2.397e-13
+ PD=7.2e-07 PS=1.49e-06
mXI42/XI519/XI88/MM1 N_XI42/NET782_XI42/XI519/XI88/MM1_d
+ N_XI42/XI519/NET104_XI42/XI519/XI88/MM1_g N_VDD_XI42/XI519/XI88/MM1_s
+ N_VDD_XI42/XI519/XI88/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13 AS=2.632e-13
+ PD=7.2e-07 PS=1.59e-06
mXI42/XI519/XI89/MM0 N_XI42/NET783_XI42/XI519/XI89/MM0_d
+ N_XI42/XI519/NET114_XI42/XI519/XI89/MM0_g N_VDD_XI42/XI519/XI89/MM0_s
+ N_VDD_XI42/XI519/XI89/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13 AS=2.397e-13
+ PD=7.2e-07 PS=1.49e-06
mXI42/XI519/XI89/MM1 N_XI42/NET783_XI42/XI519/XI89/MM1_d
+ N_XI42/XI519/NET103_XI42/XI519/XI89/MM1_g N_VDD_XI42/XI519/XI89/MM1_s
+ N_VDD_XI42/XI519/XI89/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13 AS=2.632e-13
+ PD=7.2e-07 PS=1.59e-06
mXI42/XI519/XI82/MM0 N_XI42/NET784_XI42/XI519/XI82/MM0_d
+ N_XI42/XI519/NET113_XI42/XI519/XI82/MM0_g N_VDD_XI42/XI519/XI82/MM0_s
+ N_VDD_XI42/XI519/XI82/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13 AS=2.397e-13
+ PD=7.2e-07 PS=1.49e-06
mXI42/XI519/XI82/MM1 N_XI42/NET784_XI42/XI519/XI82/MM1_d
+ N_XI42/XI519/NET36_XI42/XI519/XI82/MM1_g N_VDD_XI42/XI519/XI82/MM1_s
+ N_VDD_XI42/XI519/XI82/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13 AS=2.632e-13
+ PD=7.2e-07 PS=1.59e-06
mXI42/XI519/XI83/MM0 N_XI42/NET785_XI42/XI519/XI83/MM0_d
+ N_XI42/XI519/NET113_XI42/XI519/XI83/MM0_g N_VDD_XI42/XI519/XI83/MM0_s
+ N_VDD_XI42/XI519/XI83/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13 AS=2.397e-13
+ PD=7.2e-07 PS=1.49e-06
mXI42/XI519/XI83/MM1 N_XI42/NET785_XI42/XI519/XI83/MM1_d
+ N_XI42/XI519/NET31_XI42/XI519/XI83/MM1_g N_VDD_XI42/XI519/XI83/MM1_s
+ N_VDD_XI42/XI519/XI83/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13 AS=2.632e-13
+ PD=7.2e-07 PS=1.59e-06
mXI42/XI519/XI84/MM0 N_XI42/NET786_XI42/XI519/XI84/MM0_d
+ N_XI42/XI519/NET113_XI42/XI519/XI84/MM0_g N_VDD_XI42/XI519/XI84/MM0_s
+ N_VDD_XI42/XI519/XI84/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13 AS=2.397e-13
+ PD=7.2e-07 PS=1.49e-06
mXI42/XI519/XI84/MM1 N_XI42/NET786_XI42/XI519/XI84/MM1_d
+ N_XI42/XI519/NET104_XI42/XI519/XI84/MM1_g N_VDD_XI42/XI519/XI84/MM1_s
+ N_VDD_XI42/XI519/XI84/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13 AS=2.632e-13
+ PD=7.2e-07 PS=1.59e-06
mXI42/XI519/XI85/MM0 N_XI42/NET787_XI42/XI519/XI85/MM0_d
+ N_XI42/XI519/NET113_XI42/XI519/XI85/MM0_g N_VDD_XI42/XI519/XI85/MM0_s
+ N_VDD_XI42/XI519/XI85/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13 AS=2.397e-13
+ PD=7.2e-07 PS=1.49e-06
mXI42/XI519/XI85/MM1 N_XI42/NET787_XI42/XI519/XI85/MM1_d
+ N_XI42/XI519/NET103_XI42/XI519/XI85/MM1_g N_VDD_XI42/XI519/XI85/MM1_s
+ N_VDD_XI42/XI519/XI85/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13 AS=2.632e-13
+ PD=7.2e-07 PS=1.59e-06
mXI42/XI519/XI78/MM0 N_XI42/NET788_XI42/XI519/XI78/MM0_d
+ N_XI42/XI519/NET112_XI42/XI519/XI78/MM0_g N_VDD_XI42/XI519/XI78/MM0_s
+ N_VDD_XI42/XI519/XI78/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13 AS=2.397e-13
+ PD=7.2e-07 PS=1.49e-06
mXI42/XI519/XI78/MM1 N_XI42/NET788_XI42/XI519/XI78/MM1_d
+ N_XI42/XI519/NET36_XI42/XI519/XI78/MM1_g N_VDD_XI42/XI519/XI78/MM1_s
+ N_VDD_XI42/XI519/XI78/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13 AS=2.632e-13
+ PD=7.2e-07 PS=1.59e-06
mXI42/XI519/XI79/MM0 N_XI42/NET789_XI42/XI519/XI79/MM0_d
+ N_XI42/XI519/NET112_XI42/XI519/XI79/MM0_g N_VDD_XI42/XI519/XI79/MM0_s
+ N_VDD_XI42/XI519/XI79/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13 AS=2.397e-13
+ PD=7.2e-07 PS=1.49e-06
mXI42/XI519/XI79/MM1 N_XI42/NET789_XI42/XI519/XI79/MM1_d
+ N_XI42/XI519/NET31_XI42/XI519/XI79/MM1_g N_VDD_XI42/XI519/XI79/MM1_s
+ N_VDD_XI42/XI519/XI79/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13 AS=2.632e-13
+ PD=7.2e-07 PS=1.59e-06
mXI42/XI519/XI80/MM0 N_XI42/NET790_XI42/XI519/XI80/MM0_d
+ N_XI42/XI519/NET112_XI42/XI519/XI80/MM0_g N_VDD_XI42/XI519/XI80/MM0_s
+ N_VDD_XI42/XI519/XI80/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13 AS=2.397e-13
+ PD=7.2e-07 PS=1.49e-06
mXI42/XI519/XI80/MM1 N_XI42/NET790_XI42/XI519/XI80/MM1_d
+ N_XI42/XI519/NET104_XI42/XI519/XI80/MM1_g N_VDD_XI42/XI519/XI80/MM1_s
+ N_VDD_XI42/XI519/XI80/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13 AS=2.632e-13
+ PD=7.2e-07 PS=1.59e-06
mXI42/XI519/XI81/MM0 N_XI42/NET791_XI42/XI519/XI81/MM0_d
+ N_XI42/XI519/NET112_XI42/XI519/XI81/MM0_g N_VDD_XI42/XI519/XI81/MM0_s
+ N_VDD_XI42/XI519/XI81/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13 AS=2.397e-13
+ PD=7.2e-07 PS=1.49e-06
mXI42/XI519/XI81/MM1 N_XI42/NET791_XI42/XI519/XI81/MM1_d
+ N_XI42/XI519/NET103_XI42/XI519/XI81/MM1_g N_VDD_XI42/XI519/XI81/MM1_s
+ N_VDD_XI42/XI519/XI81/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13 AS=2.632e-13
+ PD=7.2e-07 PS=1.59e-06
mXI42/XI519/XI74/MM0 N_XI42/NET792_XI42/XI519/XI74/MM0_d
+ N_XI42/XI519/NET111_XI42/XI519/XI74/MM0_g N_VDD_XI42/XI519/XI74/MM0_s
+ N_VDD_XI42/XI519/XI74/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13 AS=2.397e-13
+ PD=7.2e-07 PS=1.49e-06
mXI42/XI519/XI74/MM1 N_XI42/NET792_XI42/XI519/XI74/MM1_d
+ N_XI42/XI519/NET36_XI42/XI519/XI74/MM1_g N_VDD_XI42/XI519/XI74/MM1_s
+ N_VDD_XI42/XI519/XI74/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13 AS=2.632e-13
+ PD=7.2e-07 PS=1.59e-06
mXI42/XI519/XI75/MM0 N_XI42/NET793_XI42/XI519/XI75/MM0_d
+ N_XI42/XI519/NET111_XI42/XI519/XI75/MM0_g N_VDD_XI42/XI519/XI75/MM0_s
+ N_VDD_XI42/XI519/XI75/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13 AS=2.397e-13
+ PD=7.2e-07 PS=1.49e-06
mXI42/XI519/XI75/MM1 N_XI42/NET793_XI42/XI519/XI75/MM1_d
+ N_XI42/XI519/NET31_XI42/XI519/XI75/MM1_g N_VDD_XI42/XI519/XI75/MM1_s
+ N_VDD_XI42/XI519/XI75/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13 AS=2.632e-13
+ PD=7.2e-07 PS=1.59e-06
mXI42/XI519/XI76/MM0 N_XI42/NET794_XI42/XI519/XI76/MM0_d
+ N_XI42/XI519/NET111_XI42/XI519/XI76/MM0_g N_VDD_XI42/XI519/XI76/MM0_s
+ N_VDD_XI42/XI519/XI76/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13 AS=2.397e-13
+ PD=7.2e-07 PS=1.49e-06
mXI42/XI519/XI76/MM1 N_XI42/NET794_XI42/XI519/XI76/MM1_d
+ N_XI42/XI519/NET104_XI42/XI519/XI76/MM1_g N_VDD_XI42/XI519/XI76/MM1_s
+ N_VDD_XI42/XI519/XI76/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13 AS=2.632e-13
+ PD=7.2e-07 PS=1.59e-06
mXI42/XI519/XI77/MM0 N_XI42/NET795_XI42/XI519/XI77/MM0_d
+ N_XI42/XI519/NET111_XI42/XI519/XI77/MM0_g N_VDD_XI42/XI519/XI77/MM0_s
+ N_VDD_XI42/XI519/XI77/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13 AS=2.397e-13
+ PD=7.2e-07 PS=1.49e-06
mXI42/XI519/XI77/MM1 N_XI42/NET795_XI42/XI519/XI77/MM1_d
+ N_XI42/XI519/NET103_XI42/XI519/XI77/MM1_g N_VDD_XI42/XI519/XI77/MM1_s
+ N_VDD_XI42/XI519/XI77/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13 AS=2.632e-13
+ PD=7.2e-07 PS=1.59e-06
mXI42/XI520/XI12/MM12 N_XI42/NET801_XI42/XI520/XI12/MM12_d
+ N_NET140_XI42/XI520/XI12/MM12_g N_VDD_XI42/XI520/XI12/MM12_s
+ N_VDD_XI42/XI519/XI86/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI42/XI520/XI12/MM13 N_XI42/NET801_XI42/XI520/XI12/MM13_d
+ N_NET138_XI42/XI520/XI12/MM13_g N_VDD_XI42/XI520/XI12/MM13_s
+ N_VDD_XI42/XI519/XI86/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13
+ AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI42/XI520/XI12/MM14 N_XI42/NET801_XI42/XI520/XI12/MM14_d
+ N_NET136_XI42/XI520/XI12/MM14_g N_VDD_XI42/XI520/XI12/MM14_s
+ N_VDD_XI42/XI519/XI86/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13
+ AS=2.726e-13 PD=5.1e-07 PS=1.63e-06
mXI42/XI520/XI13/MM12 N_XI42/NET455_XI42/XI520/XI13/MM12_d
+ N_NET140_XI42/XI520/XI13/MM12_g N_VDD_XI42/XI520/XI13/MM12_s
+ N_VDD_XI42/XI520/XI13/MM12_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI42/XI520/XI13/MM13 N_XI42/NET455_XI42/XI520/XI13/MM13_d
+ N_NET138_XI42/XI520/XI13/MM13_g N_VDD_XI42/XI520/XI13/MM13_s
+ N_VDD_XI42/XI520/XI13/MM12_b P_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13
+ AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI42/XI520/XI13/MM14 N_XI42/NET455_XI42/XI520/XI13/MM14_d
+ N_NET135_XI42/XI520/XI13/MM14_g N_VDD_XI42/XI520/XI13/MM14_s
+ N_VDD_XI42/XI520/XI13/MM12_b P_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13
+ AS=2.726e-13 PD=5.1e-07 PS=1.63e-06
mXI42/XI520/XI14/MM12 N_XI42/NET803_XI42/XI520/XI14/MM12_d
+ N_NET140_XI42/XI520/XI14/MM12_g N_VDD_XI42/XI520/XI14/MM12_s
+ N_VDD_XI42/XI520/XI14/MM12_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI42/XI520/XI14/MM13 N_XI42/NET803_XI42/XI520/XI14/MM13_d
+ N_NET137_XI42/XI520/XI14/MM13_g N_VDD_XI42/XI520/XI14/MM13_s
+ N_VDD_XI42/XI520/XI14/MM12_b P_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13
+ AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI42/XI520/XI14/MM14 N_XI42/NET803_XI42/XI520/XI14/MM14_d
+ N_NET136_XI42/XI520/XI14/MM14_g N_VDD_XI42/XI520/XI14/MM14_s
+ N_VDD_XI42/XI520/XI14/MM12_b P_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13
+ AS=2.726e-13 PD=5.1e-07 PS=1.63e-06
mXI42/XI520/XI15/MM12 N_XI42/NET245_XI42/XI520/XI15/MM12_d
+ N_NET140_XI42/XI520/XI15/MM12_g N_VDD_XI42/XI520/XI15/MM12_s
+ N_VDD_XI42/XI520/XI14/MM12_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI42/XI520/XI15/MM13 N_XI42/NET245_XI42/XI520/XI15/MM13_d
+ N_NET137_XI42/XI520/XI15/MM13_g N_VDD_XI42/XI520/XI15/MM13_s
+ N_VDD_XI42/XI520/XI14/MM12_b P_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13
+ AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI42/XI520/XI15/MM14 N_XI42/NET245_XI42/XI520/XI15/MM14_d
+ N_NET135_XI42/XI520/XI15/MM14_g N_VDD_XI42/XI520/XI15/MM14_s
+ N_VDD_XI42/XI520/XI14/MM12_b P_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13
+ AS=2.726e-13 PD=5.1e-07 PS=1.63e-06
mXI42/XI520/XI16/MM12 N_XI42/NET802_XI42/XI520/XI16/MM12_d
+ N_NET139_XI42/XI520/XI16/MM12_g N_VDD_XI42/XI520/XI16/MM12_s
+ N_VDD_XI42/XI520/XI16/MM12_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI42/XI520/XI16/MM13 N_XI42/NET802_XI42/XI520/XI16/MM13_d
+ N_NET138_XI42/XI520/XI16/MM13_g N_VDD_XI42/XI520/XI16/MM13_s
+ N_VDD_XI42/XI520/XI16/MM12_b P_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13
+ AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI42/XI520/XI16/MM14 N_XI42/NET802_XI42/XI520/XI16/MM14_d
+ N_NET136_XI42/XI520/XI16/MM14_g N_VDD_XI42/XI520/XI16/MM14_s
+ N_VDD_XI42/XI520/XI16/MM12_b P_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13
+ AS=2.726e-13 PD=5.1e-07 PS=1.63e-06
mXI42/XI520/XI17/MM12 N_XI42/NET375_XI42/XI520/XI17/MM12_d
+ N_NET139_XI42/XI520/XI17/MM12_g N_VDD_XI42/XI520/XI17/MM12_s
+ N_VDD_XI42/XI520/XI16/MM12_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI42/XI520/XI17/MM13 N_XI42/NET375_XI42/XI520/XI17/MM13_d
+ N_NET138_XI42/XI520/XI17/MM13_g N_VDD_XI42/XI520/XI17/MM13_s
+ N_VDD_XI42/XI520/XI16/MM12_b P_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13
+ AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI42/XI520/XI17/MM14 N_XI42/NET375_XI42/XI520/XI17/MM14_d
+ N_NET135_XI42/XI520/XI17/MM14_g N_VDD_XI42/XI520/XI17/MM14_s
+ N_VDD_XI42/XI520/XI16/MM12_b P_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13
+ AS=2.726e-13 PD=5.1e-07 PS=1.63e-06
mXI42/XI520/XI18/MM12 N_XI42/NET535_XI42/XI520/XI18/MM12_d
+ N_NET139_XI42/XI520/XI18/MM12_g N_VDD_XI42/XI520/XI18/MM12_s
+ N_VDD_XI42/XI520/XI18/MM12_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI42/XI520/XI18/MM13 N_XI42/NET535_XI42/XI520/XI18/MM13_d
+ N_NET137_XI42/XI520/XI18/MM13_g N_VDD_XI42/XI520/XI18/MM13_s
+ N_VDD_XI42/XI520/XI18/MM12_b P_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13
+ AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI42/XI520/XI18/MM14 N_XI42/NET535_XI42/XI520/XI18/MM14_d
+ N_NET136_XI42/XI520/XI18/MM14_g N_VDD_XI42/XI520/XI18/MM14_s
+ N_VDD_XI42/XI520/XI18/MM12_b P_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13
+ AS=2.726e-13 PD=5.1e-07 PS=1.63e-06
mXI42/XI520/XI19/MM12 N_XI42/NET180_XI42/XI520/XI19/MM12_d
+ N_NET139_XI42/XI520/XI19/MM12_g N_VDD_XI42/XI520/XI19/MM12_s
+ N_VDD_XI42/XI520/XI18/MM12_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI42/XI520/XI19/MM13 N_XI42/NET180_XI42/XI520/XI19/MM13_d
+ N_NET137_XI42/XI520/XI19/MM13_g N_VDD_XI42/XI520/XI19/MM13_s
+ N_VDD_XI42/XI520/XI18/MM12_b P_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13
+ AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI42/XI520/XI19/MM14 N_XI42/NET180_XI42/XI520/XI19/MM14_d
+ N_NET135_XI42/XI520/XI19/MM14_g N_VDD_XI42/XI520/XI19/MM14_s
+ N_VDD_XI42/XI520/XI18/MM12_b P_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13
+ AS=2.726e-13 PD=5.1e-07 PS=1.63e-06
mXI54/XI0/XI8/XI3/MM1 N_XI54/XI0/XI8/NET12_XI54/XI0/XI8/XI3/MM1_d
+ N_XI54/XI0/NET2_XI54/XI0/XI8/XI3/MM1_g N_VDD_XI54/XI0/XI8/XI3/MM1_s
+ N_VDD_XI30/XI67/MM2_b P_18 L=1.8e-07 W=4.7e-07 AD=1.68025e-13 AS=2.303e-13
+ PD=7.15e-07 PS=1.45e-06
mXI54/XI0/XI7/XI3/MM1 N_XI54/XI0/XI7/NET12_XI54/XI0/XI7/XI3/MM1_d
+ N_NET062_XI54/XI0/XI7/XI3/MM1_g N_VDD_XI54/XI0/XI7/XI3/MM1_s
+ N_VDD_XI30/XI67/MM2_b P_18 L=1.8e-07 W=4.7e-07 AD=1.68025e-13 AS=2.5145e-13
+ PD=7.15e-07 PS=1.54e-06
mXI54/XI0/XI6/MM0 N_XI54/XI0/NET2_XI54/XI0/XI6/MM0_d N_NET062_XI54/XI0/XI6/MM0_g
+ N_VDD_XI54/XI0/XI6/MM0_s N_VDD_XI30/XI67/MM2_b P_18 L=1.8e-07 W=1.85e-06
+ AD=9.435e-13 AS=9.435e-13 PD=2.87e-06 PS=2.87e-06
mXI42/XI649/XI2/MM0 N_XI42/NET0373_XI42/XI649/XI2/MM0_d
+ N_NET070_XI42/XI649/XI2/MM0_g N_VDD_XI42/XI649/XI2/MM0_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13 AS=2.397e-13
+ PD=7.2e-07 PS=1.49e-06
mXI42/XI649/XI2/MM1 N_XI42/NET0373_XI42/XI649/XI2/MM1_d
+ N_XI42/NET0388_XI42/XI649/XI2/MM1_g N_VDD_XI42/XI649/XI2/MM1_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=1.692e-13 AS=2.632e-13
+ PD=7.2e-07 PS=1.59e-06
mXI57/XI0/MM3 N_XI57/NET19_XI57/XI0/MM3_d N_NET068_XI57/XI0/MM3_g
+ N_VDD_XI57/XI0/MM3_s N_VDD_XI30/XI67/MM2_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.35e-13 AS=1.7625e-13 PD=1.47e-06 PS=7.5e-07
mXI57/XI0/MM2 N_XI57/NET19_XI57/XI0/MM2_d N_NET062_XI57/XI0/MM2_g
+ N_VDD_XI57/XI0/MM2_s N_VDD_XI30/XI67/MM2_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.3735e-13 AS=1.7625e-13 PD=1.48e-06 PS=7.5e-07
mXI57/XI0/MM1 N_NET062_XI57/XI0/MM1_d N_XI57/NET19_XI57/XI0/MM1_g
+ N_VDD_XI57/XI0/MM1_s N_VDD_XI30/XI67/MM2_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.3735e-13 AS=1.7625e-13 PD=1.48e-06 PS=7.5e-07
mXI57/XI0/MM0 N_NET062_XI57/XI0/MM0_d N_NET068_XI57/XI0/MM0_g
+ N_VDD_XI57/XI0/MM0_s N_VDD_XI30/XI67/MM2_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.35e-13 AS=1.7625e-13 PD=1.47e-06 PS=7.5e-07
mXI42/XI649/XI3/MM0 N_NET0390_XI42/XI649/XI3/MM0_d
+ N_XI42/NET0373_XI42/XI649/XI3/MM0_g N_VDD_XI42/XI649/XI3/MM0_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=1.85e-06 AD=9.435e-13 AS=9.435e-13
+ PD=2.87e-06 PS=2.87e-06
mXI42/XI648/MM7 N_XI42/XI648/NET21_XI42/XI648/MM7_d
+ N_XI42/NET780_XI42/XI648/MM7_g N_VDD_XI42/XI648/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI584/MM7 N_XI42/XI584/NET21_XI42/XI584/MM7_d
+ N_XI42/NET780_XI42/XI584/MM7_g N_VDD_XI42/XI584/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI616/MM7 N_XI42/XI616/NET21_XI42/XI616/MM7_d
+ N_XI42/NET780_XI42/XI616/MM7_g N_VDD_XI42/XI616/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI552/MM7 N_XI42/XI552/NET21_XI42/XI552/MM7_d
+ N_XI42/NET780_XI42/XI552/MM7_g N_VDD_XI42/XI552/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI632/MM7 N_XI42/XI632/NET21_XI42/XI632/MM7_d
+ N_XI42/NET780_XI42/XI632/MM7_g N_VDD_XI42/XI632/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI568/MM7 N_XI42/XI568/NET21_XI42/XI568/MM7_d
+ N_XI42/NET780_XI42/XI568/MM7_g N_VDD_XI42/XI568/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI600/MM7 N_XI42/XI600/NET21_XI42/XI600/MM7_d
+ N_XI42/NET780_XI42/XI600/MM7_g N_VDD_XI42/XI600/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI536/MM7 N_XI42/XI536/NET21_XI42/XI536/MM7_d
+ N_XI42/NET780_XI42/XI536/MM7_g N_VDD_XI42/XI536/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI647/MM7 N_XI42/XI647/NET21_XI42/XI647/MM7_d
+ N_XI42/NET781_XI42/XI647/MM7_g N_VDD_XI42/XI647/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI583/MM7 N_XI42/XI583/NET21_XI42/XI583/MM7_d
+ N_XI42/NET781_XI42/XI583/MM7_g N_VDD_XI42/XI583/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI615/MM7 N_XI42/XI615/NET21_XI42/XI615/MM7_d
+ N_XI42/NET781_XI42/XI615/MM7_g N_VDD_XI42/XI615/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI551/MM7 N_XI42/XI551/NET21_XI42/XI551/MM7_d
+ N_XI42/NET781_XI42/XI551/MM7_g N_VDD_XI42/XI551/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI631/MM7 N_XI42/XI631/NET21_XI42/XI631/MM7_d
+ N_XI42/NET781_XI42/XI631/MM7_g N_VDD_XI42/XI631/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI567/MM7 N_XI42/XI567/NET21_XI42/XI567/MM7_d
+ N_XI42/NET781_XI42/XI567/MM7_g N_VDD_XI42/XI567/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI599/MM7 N_XI42/XI599/NET21_XI42/XI599/MM7_d
+ N_XI42/NET781_XI42/XI599/MM7_g N_VDD_XI42/XI599/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI535/MM7 N_XI42/XI535/NET21_XI42/XI535/MM7_d
+ N_XI42/NET781_XI42/XI535/MM7_g N_VDD_XI42/XI535/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI646/MM7 N_XI42/XI646/NET21_XI42/XI646/MM7_d
+ N_XI42/NET782_XI42/XI646/MM7_g N_VDD_XI42/XI646/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI582/MM7 N_XI42/XI582/NET21_XI42/XI582/MM7_d
+ N_XI42/NET782_XI42/XI582/MM7_g N_VDD_XI42/XI582/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI614/MM7 N_XI42/XI614/NET21_XI42/XI614/MM7_d
+ N_XI42/NET782_XI42/XI614/MM7_g N_VDD_XI42/XI614/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI550/MM7 N_XI42/XI550/NET21_XI42/XI550/MM7_d
+ N_XI42/NET782_XI42/XI550/MM7_g N_VDD_XI42/XI550/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI630/MM7 N_XI42/XI630/NET21_XI42/XI630/MM7_d
+ N_XI42/NET782_XI42/XI630/MM7_g N_VDD_XI42/XI630/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI566/MM7 N_XI42/XI566/NET21_XI42/XI566/MM7_d
+ N_XI42/NET782_XI42/XI566/MM7_g N_VDD_XI42/XI566/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI598/MM7 N_XI42/XI598/NET21_XI42/XI598/MM7_d
+ N_XI42/NET782_XI42/XI598/MM7_g N_VDD_XI42/XI598/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI534/MM7 N_XI42/XI534/NET21_XI42/XI534/MM7_d
+ N_XI42/NET782_XI42/XI534/MM7_g N_VDD_XI42/XI534/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI645/MM7 N_XI42/XI645/NET21_XI42/XI645/MM7_d
+ N_XI42/NET783_XI42/XI645/MM7_g N_VDD_XI42/XI645/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI581/MM7 N_XI42/XI581/NET21_XI42/XI581/MM7_d
+ N_XI42/NET783_XI42/XI581/MM7_g N_VDD_XI42/XI581/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI613/MM7 N_XI42/XI613/NET21_XI42/XI613/MM7_d
+ N_XI42/NET783_XI42/XI613/MM7_g N_VDD_XI42/XI613/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI549/MM7 N_XI42/XI549/NET21_XI42/XI549/MM7_d
+ N_XI42/NET783_XI42/XI549/MM7_g N_VDD_XI42/XI549/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI629/MM7 N_XI42/XI629/NET21_XI42/XI629/MM7_d
+ N_XI42/NET783_XI42/XI629/MM7_g N_VDD_XI42/XI629/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI565/MM7 N_XI42/XI565/NET21_XI42/XI565/MM7_d
+ N_XI42/NET783_XI42/XI565/MM7_g N_VDD_XI42/XI565/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI597/MM7 N_XI42/XI597/NET21_XI42/XI597/MM7_d
+ N_XI42/NET783_XI42/XI597/MM7_g N_VDD_XI42/XI597/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI533/MM7 N_XI42/XI533/NET21_XI42/XI533/MM7_d
+ N_XI42/NET783_XI42/XI533/MM7_g N_VDD_XI42/XI533/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI644/MM7 N_XI42/XI644/NET21_XI42/XI644/MM7_d
+ N_XI42/NET784_XI42/XI644/MM7_g N_VDD_XI42/XI644/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI580/MM7 N_XI42/XI580/NET21_XI42/XI580/MM7_d
+ N_XI42/NET784_XI42/XI580/MM7_g N_VDD_XI42/XI580/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI612/MM7 N_XI42/XI612/NET21_XI42/XI612/MM7_d
+ N_XI42/NET784_XI42/XI612/MM7_g N_VDD_XI42/XI612/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI548/MM7 N_XI42/XI548/NET21_XI42/XI548/MM7_d
+ N_XI42/NET784_XI42/XI548/MM7_g N_VDD_XI42/XI548/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI628/MM7 N_XI42/XI628/NET21_XI42/XI628/MM7_d
+ N_XI42/NET784_XI42/XI628/MM7_g N_VDD_XI42/XI628/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI564/MM7 N_XI42/XI564/NET21_XI42/XI564/MM7_d
+ N_XI42/NET784_XI42/XI564/MM7_g N_VDD_XI42/XI564/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI596/MM7 N_XI42/XI596/NET21_XI42/XI596/MM7_d
+ N_XI42/NET784_XI42/XI596/MM7_g N_VDD_XI42/XI596/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI532/MM7 N_XI42/XI532/NET21_XI42/XI532/MM7_d
+ N_XI42/NET784_XI42/XI532/MM7_g N_VDD_XI42/XI532/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI643/MM7 N_XI42/XI643/NET21_XI42/XI643/MM7_d
+ N_XI42/NET785_XI42/XI643/MM7_g N_VDD_XI42/XI643/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI579/MM7 N_XI42/XI579/NET21_XI42/XI579/MM7_d
+ N_XI42/NET785_XI42/XI579/MM7_g N_VDD_XI42/XI579/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI611/MM7 N_XI42/XI611/NET21_XI42/XI611/MM7_d
+ N_XI42/NET785_XI42/XI611/MM7_g N_VDD_XI42/XI611/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI547/MM7 N_XI42/XI547/NET21_XI42/XI547/MM7_d
+ N_XI42/NET785_XI42/XI547/MM7_g N_VDD_XI42/XI547/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI627/MM7 N_XI42/XI627/NET21_XI42/XI627/MM7_d
+ N_XI42/NET785_XI42/XI627/MM7_g N_VDD_XI42/XI627/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI563/MM7 N_XI42/XI563/NET21_XI42/XI563/MM7_d
+ N_XI42/NET785_XI42/XI563/MM7_g N_VDD_XI42/XI563/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI595/MM7 N_XI42/XI595/NET21_XI42/XI595/MM7_d
+ N_XI42/NET785_XI42/XI595/MM7_g N_VDD_XI42/XI595/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI531/MM7 N_XI42/XI531/NET21_XI42/XI531/MM7_d
+ N_XI42/NET785_XI42/XI531/MM7_g N_VDD_XI42/XI531/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI642/MM7 N_XI42/XI642/NET21_XI42/XI642/MM7_d
+ N_XI42/NET786_XI42/XI642/MM7_g N_VDD_XI42/XI642/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI578/MM7 N_XI42/XI578/NET21_XI42/XI578/MM7_d
+ N_XI42/NET786_XI42/XI578/MM7_g N_VDD_XI42/XI578/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI610/MM7 N_XI42/XI610/NET21_XI42/XI610/MM7_d
+ N_XI42/NET786_XI42/XI610/MM7_g N_VDD_XI42/XI610/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI546/MM7 N_XI42/XI546/NET21_XI42/XI546/MM7_d
+ N_XI42/NET786_XI42/XI546/MM7_g N_VDD_XI42/XI546/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI626/MM7 N_XI42/XI626/NET21_XI42/XI626/MM7_d
+ N_XI42/NET786_XI42/XI626/MM7_g N_VDD_XI42/XI626/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI562/MM7 N_XI42/XI562/NET21_XI42/XI562/MM7_d
+ N_XI42/NET786_XI42/XI562/MM7_g N_VDD_XI42/XI562/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI594/MM7 N_XI42/XI594/NET21_XI42/XI594/MM7_d
+ N_XI42/NET786_XI42/XI594/MM7_g N_VDD_XI42/XI594/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI530/MM7 N_XI42/XI530/NET21_XI42/XI530/MM7_d
+ N_XI42/NET786_XI42/XI530/MM7_g N_VDD_XI42/XI530/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI641/MM7 N_XI42/XI641/NET21_XI42/XI641/MM7_d
+ N_XI42/NET787_XI42/XI641/MM7_g N_VDD_XI42/XI641/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI577/MM7 N_XI42/XI577/NET21_XI42/XI577/MM7_d
+ N_XI42/NET787_XI42/XI577/MM7_g N_VDD_XI42/XI577/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI609/MM7 N_XI42/XI609/NET21_XI42/XI609/MM7_d
+ N_XI42/NET787_XI42/XI609/MM7_g N_VDD_XI42/XI609/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI545/MM7 N_XI42/XI545/NET21_XI42/XI545/MM7_d
+ N_XI42/NET787_XI42/XI545/MM7_g N_VDD_XI42/XI545/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI625/MM7 N_XI42/XI625/NET21_XI42/XI625/MM7_d
+ N_XI42/NET787_XI42/XI625/MM7_g N_VDD_XI42/XI625/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI561/MM7 N_XI42/XI561/NET21_XI42/XI561/MM7_d
+ N_XI42/NET787_XI42/XI561/MM7_g N_VDD_XI42/XI561/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI593/MM7 N_XI42/XI593/NET21_XI42/XI593/MM7_d
+ N_XI42/NET787_XI42/XI593/MM7_g N_VDD_XI42/XI593/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI529/MM7 N_XI42/XI529/NET21_XI42/XI529/MM7_d
+ N_XI42/NET787_XI42/XI529/MM7_g N_VDD_XI42/XI529/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI640/MM7 N_XI42/XI640/NET21_XI42/XI640/MM7_d
+ N_XI42/NET788_XI42/XI640/MM7_g N_VDD_XI42/XI640/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI576/MM7 N_XI42/XI576/NET21_XI42/XI576/MM7_d
+ N_XI42/NET788_XI42/XI576/MM7_g N_VDD_XI42/XI576/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI608/MM7 N_XI42/XI608/NET21_XI42/XI608/MM7_d
+ N_XI42/NET788_XI42/XI608/MM7_g N_VDD_XI42/XI608/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI544/MM7 N_XI42/XI544/NET21_XI42/XI544/MM7_d
+ N_XI42/NET788_XI42/XI544/MM7_g N_VDD_XI42/XI544/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI624/MM7 N_XI42/XI624/NET21_XI42/XI624/MM7_d
+ N_XI42/NET788_XI42/XI624/MM7_g N_VDD_XI42/XI624/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI560/MM7 N_XI42/XI560/NET21_XI42/XI560/MM7_d
+ N_XI42/NET788_XI42/XI560/MM7_g N_VDD_XI42/XI560/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI592/MM7 N_XI42/XI592/NET21_XI42/XI592/MM7_d
+ N_XI42/NET788_XI42/XI592/MM7_g N_VDD_XI42/XI592/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI528/MM7 N_XI42/XI528/NET21_XI42/XI528/MM7_d
+ N_XI42/NET788_XI42/XI528/MM7_g N_VDD_XI42/XI528/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI639/MM7 N_XI42/XI639/NET21_XI42/XI639/MM7_d
+ N_XI42/NET789_XI42/XI639/MM7_g N_VDD_XI42/XI639/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI575/MM7 N_XI42/XI575/NET21_XI42/XI575/MM7_d
+ N_XI42/NET789_XI42/XI575/MM7_g N_VDD_XI42/XI575/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI607/MM7 N_XI42/XI607/NET21_XI42/XI607/MM7_d
+ N_XI42/NET789_XI42/XI607/MM7_g N_VDD_XI42/XI607/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI543/MM7 N_XI42/XI543/NET21_XI42/XI543/MM7_d
+ N_XI42/NET789_XI42/XI543/MM7_g N_VDD_XI42/XI543/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI623/MM7 N_XI42/XI623/NET21_XI42/XI623/MM7_d
+ N_XI42/NET789_XI42/XI623/MM7_g N_VDD_XI42/XI623/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI559/MM7 N_XI42/XI559/NET21_XI42/XI559/MM7_d
+ N_XI42/NET789_XI42/XI559/MM7_g N_VDD_XI42/XI559/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI591/MM7 N_XI42/XI591/NET21_XI42/XI591/MM7_d
+ N_XI42/NET789_XI42/XI591/MM7_g N_VDD_XI42/XI591/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI527/MM7 N_XI42/XI527/NET21_XI42/XI527/MM7_d
+ N_XI42/NET789_XI42/XI527/MM7_g N_VDD_XI42/XI527/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI638/MM7 N_XI42/XI638/NET21_XI42/XI638/MM7_d
+ N_XI42/NET790_XI42/XI638/MM7_g N_VDD_XI42/XI638/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI574/MM7 N_XI42/XI574/NET21_XI42/XI574/MM7_d
+ N_XI42/NET790_XI42/XI574/MM7_g N_VDD_XI42/XI574/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI606/MM7 N_XI42/XI606/NET21_XI42/XI606/MM7_d
+ N_XI42/NET790_XI42/XI606/MM7_g N_VDD_XI42/XI606/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI542/MM7 N_XI42/XI542/NET21_XI42/XI542/MM7_d
+ N_XI42/NET790_XI42/XI542/MM7_g N_VDD_XI42/XI542/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI622/MM7 N_XI42/XI622/NET21_XI42/XI622/MM7_d
+ N_XI42/NET790_XI42/XI622/MM7_g N_VDD_XI42/XI622/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI558/MM7 N_XI42/XI558/NET21_XI42/XI558/MM7_d
+ N_XI42/NET790_XI42/XI558/MM7_g N_VDD_XI42/XI558/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI590/MM7 N_XI42/XI590/NET21_XI42/XI590/MM7_d
+ N_XI42/NET790_XI42/XI590/MM7_g N_VDD_XI42/XI590/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI526/MM7 N_XI42/XI526/NET21_XI42/XI526/MM7_d
+ N_XI42/NET790_XI42/XI526/MM7_g N_VDD_XI42/XI526/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI637/MM7 N_XI42/XI637/NET21_XI42/XI637/MM7_d
+ N_XI42/NET791_XI42/XI637/MM7_g N_VDD_XI42/XI637/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI573/MM7 N_XI42/XI573/NET21_XI42/XI573/MM7_d
+ N_XI42/NET791_XI42/XI573/MM7_g N_VDD_XI42/XI573/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI605/MM7 N_XI42/XI605/NET21_XI42/XI605/MM7_d
+ N_XI42/NET791_XI42/XI605/MM7_g N_VDD_XI42/XI605/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI541/MM7 N_XI42/XI541/NET21_XI42/XI541/MM7_d
+ N_XI42/NET791_XI42/XI541/MM7_g N_VDD_XI42/XI541/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI621/MM7 N_XI42/XI621/NET21_XI42/XI621/MM7_d
+ N_XI42/NET791_XI42/XI621/MM7_g N_VDD_XI42/XI621/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI557/MM7 N_XI42/XI557/NET21_XI42/XI557/MM7_d
+ N_XI42/NET791_XI42/XI557/MM7_g N_VDD_XI42/XI557/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI589/MM7 N_XI42/XI589/NET21_XI42/XI589/MM7_d
+ N_XI42/NET791_XI42/XI589/MM7_g N_VDD_XI42/XI589/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI525/MM7 N_XI42/XI525/NET21_XI42/XI525/MM7_d
+ N_XI42/NET791_XI42/XI525/MM7_g N_VDD_XI42/XI525/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI636/MM7 N_XI42/XI636/NET21_XI42/XI636/MM7_d
+ N_XI42/NET792_XI42/XI636/MM7_g N_VDD_XI42/XI636/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI572/MM7 N_XI42/XI572/NET21_XI42/XI572/MM7_d
+ N_XI42/NET792_XI42/XI572/MM7_g N_VDD_XI42/XI572/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI604/MM7 N_XI42/XI604/NET21_XI42/XI604/MM7_d
+ N_XI42/NET792_XI42/XI604/MM7_g N_VDD_XI42/XI604/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI540/MM7 N_XI42/XI540/NET21_XI42/XI540/MM7_d
+ N_XI42/NET792_XI42/XI540/MM7_g N_VDD_XI42/XI540/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI620/MM7 N_XI42/XI620/NET21_XI42/XI620/MM7_d
+ N_XI42/NET792_XI42/XI620/MM7_g N_VDD_XI42/XI620/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI556/MM7 N_XI42/XI556/NET21_XI42/XI556/MM7_d
+ N_XI42/NET792_XI42/XI556/MM7_g N_VDD_XI42/XI556/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI588/MM7 N_XI42/XI588/NET21_XI42/XI588/MM7_d
+ N_XI42/NET792_XI42/XI588/MM7_g N_VDD_XI42/XI588/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI524/MM7 N_XI42/XI524/NET21_XI42/XI524/MM7_d
+ N_XI42/NET792_XI42/XI524/MM7_g N_VDD_XI42/XI524/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI635/MM7 N_XI42/XI635/NET21_XI42/XI635/MM7_d
+ N_XI42/NET793_XI42/XI635/MM7_g N_VDD_XI42/XI635/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI571/MM7 N_XI42/XI571/NET21_XI42/XI571/MM7_d
+ N_XI42/NET793_XI42/XI571/MM7_g N_VDD_XI42/XI571/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI603/MM7 N_XI42/XI603/NET21_XI42/XI603/MM7_d
+ N_XI42/NET793_XI42/XI603/MM7_g N_VDD_XI42/XI603/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI539/MM7 N_XI42/XI539/NET21_XI42/XI539/MM7_d
+ N_XI42/NET793_XI42/XI539/MM7_g N_VDD_XI42/XI539/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI619/MM7 N_XI42/XI619/NET21_XI42/XI619/MM7_d
+ N_XI42/NET793_XI42/XI619/MM7_g N_VDD_XI42/XI619/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI555/MM7 N_XI42/XI555/NET21_XI42/XI555/MM7_d
+ N_XI42/NET793_XI42/XI555/MM7_g N_VDD_XI42/XI555/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI587/MM7 N_XI42/XI587/NET21_XI42/XI587/MM7_d
+ N_XI42/NET793_XI42/XI587/MM7_g N_VDD_XI42/XI587/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI523/MM7 N_XI42/XI523/NET21_XI42/XI523/MM7_d
+ N_XI42/NET793_XI42/XI523/MM7_g N_VDD_XI42/XI523/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI634/MM7 N_XI42/XI634/NET21_XI42/XI634/MM7_d
+ N_XI42/NET794_XI42/XI634/MM7_g N_VDD_XI42/XI634/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI570/MM7 N_XI42/XI570/NET21_XI42/XI570/MM7_d
+ N_XI42/NET794_XI42/XI570/MM7_g N_VDD_XI42/XI570/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI602/MM7 N_XI42/XI602/NET21_XI42/XI602/MM7_d
+ N_XI42/NET794_XI42/XI602/MM7_g N_VDD_XI42/XI602/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI538/MM7 N_XI42/XI538/NET21_XI42/XI538/MM7_d
+ N_XI42/NET794_XI42/XI538/MM7_g N_VDD_XI42/XI538/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI618/MM7 N_XI42/XI618/NET21_XI42/XI618/MM7_d
+ N_XI42/NET794_XI42/XI618/MM7_g N_VDD_XI42/XI618/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI554/MM7 N_XI42/XI554/NET21_XI42/XI554/MM7_d
+ N_XI42/NET794_XI42/XI554/MM7_g N_VDD_XI42/XI554/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI586/MM7 N_XI42/XI586/NET21_XI42/XI586/MM7_d
+ N_XI42/NET794_XI42/XI586/MM7_g N_VDD_XI42/XI586/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI522/MM7 N_XI42/XI522/NET21_XI42/XI522/MM7_d
+ N_XI42/NET794_XI42/XI522/MM7_g N_VDD_XI42/XI522/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI633/MM7 N_XI42/XI633/NET21_XI42/XI633/MM7_d
+ N_XI42/NET795_XI42/XI633/MM7_g N_VDD_XI42/XI633/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI569/MM7 N_XI42/XI569/NET21_XI42/XI569/MM7_d
+ N_XI42/NET795_XI42/XI569/MM7_g N_VDD_XI42/XI569/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI601/MM7 N_XI42/XI601/NET21_XI42/XI601/MM7_d
+ N_XI42/NET795_XI42/XI601/MM7_g N_VDD_XI42/XI601/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI537/MM7 N_XI42/XI537/NET21_XI42/XI537/MM7_d
+ N_XI42/NET795_XI42/XI537/MM7_g N_VDD_XI42/XI537/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI617/MM7 N_XI42/XI617/NET21_XI42/XI617/MM7_d
+ N_XI42/NET795_XI42/XI617/MM7_g N_VDD_XI42/XI617/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI553/MM7 N_XI42/XI553/NET21_XI42/XI553/MM7_d
+ N_XI42/NET795_XI42/XI553/MM7_g N_VDD_XI42/XI553/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI585/MM7 N_XI42/XI585/NET21_XI42/XI585/MM7_d
+ N_XI42/NET795_XI42/XI585/MM7_g N_VDD_XI42/XI585/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI521/MM7 N_XI42/XI521/NET21_XI42/XI521/MM7_d
+ N_XI42/NET795_XI42/XI521/MM7_g N_VDD_XI42/XI521/MM7_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=7.05e-14 AS=2.632e-13
+ PD=3e-07 PS=1.59e-06
mXI42/XI648/MM6 N_XI42/NET01023_XI42/XI648/MM6_d N_XI42/NET801_XI42/XI648/MM6_g
+ N_XI42/XI648/NET21_XI42/XI648/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI584/MM6 N_NET280_XI42/XI584/MM6_d N_XI42/NET455_XI42/XI584/MM6_g
+ N_XI42/XI584/NET21_XI42/XI584/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI616/MM6 N_NET281_XI42/XI616/MM6_d N_XI42/NET803_XI42/XI616/MM6_g
+ N_XI42/XI616/NET21_XI42/XI616/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI552/MM6 N_NET282_XI42/XI552/MM6_d N_XI42/NET245_XI42/XI552/MM6_g
+ N_XI42/XI552/NET21_XI42/XI552/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI632/MM6 N_NET153_XI42/XI632/MM6_d N_XI42/NET802_XI42/XI632/MM6_g
+ N_XI42/XI632/NET21_XI42/XI632/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI568/MM6 N_NET284_XI42/XI568/MM6_d N_XI42/NET375_XI42/XI568/MM6_g
+ N_XI42/XI568/NET21_XI42/XI568/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI600/MM6 N_NET285_XI42/XI600/MM6_d N_XI42/NET535_XI42/XI600/MM6_g
+ N_XI42/XI600/NET21_XI42/XI600/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI536/MM6 N_NET286_XI42/XI536/MM6_d N_XI42/NET180_XI42/XI536/MM6_g
+ N_XI42/XI536/NET21_XI42/XI536/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI647/MM6 N_NET287_XI42/XI647/MM6_d N_XI42/NET801_XI42/XI647/MM6_g
+ N_XI42/XI647/NET21_XI42/XI647/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI583/MM6 N_NET158_XI42/XI583/MM6_d N_XI42/NET455_XI42/XI583/MM6_g
+ N_XI42/XI583/NET21_XI42/XI583/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI615/MM6 N_NET159_XI42/XI615/MM6_d N_XI42/NET803_XI42/XI615/MM6_g
+ N_XI42/XI615/NET21_XI42/XI615/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI551/MM6 N_NET160_XI42/XI551/MM6_d N_XI42/NET245_XI42/XI551/MM6_g
+ N_XI42/XI551/NET21_XI42/XI551/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI631/MM6 N_NET291_XI42/XI631/MM6_d N_XI42/NET802_XI42/XI631/MM6_g
+ N_XI42/XI631/NET21_XI42/XI631/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI567/MM6 N_NET162_XI42/XI567/MM6_d N_XI42/NET375_XI42/XI567/MM6_g
+ N_XI42/XI567/NET21_XI42/XI567/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI599/MM6 N_NET293_XI42/XI599/MM6_d N_XI42/NET535_XI42/XI599/MM6_g
+ N_XI42/XI599/NET21_XI42/XI599/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI535/MM6 N_NET294_XI42/XI535/MM6_d N_XI42/NET180_XI42/XI535/MM6_g
+ N_XI42/XI535/NET21_XI42/XI535/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI646/MM6 N_NET295_XI42/XI646/MM6_d N_XI42/NET801_XI42/XI646/MM6_g
+ N_XI42/XI646/NET21_XI42/XI646/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI582/MM6 N_NET296_XI42/XI582/MM6_d N_XI42/NET455_XI42/XI582/MM6_g
+ N_XI42/XI582/NET21_XI42/XI582/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI614/MM6 N_NET297_XI42/XI614/MM6_d N_XI42/NET803_XI42/XI614/MM6_g
+ N_XI42/XI614/NET21_XI42/XI614/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI550/MM6 N_NET298_XI42/XI550/MM6_d N_XI42/NET245_XI42/XI550/MM6_g
+ N_XI42/XI550/NET21_XI42/XI550/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI630/MM6 N_NET299_XI42/XI630/MM6_d N_XI42/NET802_XI42/XI630/MM6_g
+ N_XI42/XI630/NET21_XI42/XI630/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI566/MM6 N_NET170_XI42/XI566/MM6_d N_XI42/NET375_XI42/XI566/MM6_g
+ N_XI42/XI566/NET21_XI42/XI566/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI598/MM6 N_NET171_XI42/XI598/MM6_d N_XI42/NET535_XI42/XI598/MM6_g
+ N_XI42/XI598/NET21_XI42/XI598/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI534/MM6 N_NET172_XI42/XI534/MM6_d N_XI42/NET180_XI42/XI534/MM6_g
+ N_XI42/XI534/NET21_XI42/XI534/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI645/MM6 N_NET303_XI42/XI645/MM6_d N_XI42/NET801_XI42/XI645/MM6_g
+ N_XI42/XI645/NET21_XI42/XI645/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI581/MM6 N_NET304_XI42/XI581/MM6_d N_XI42/NET455_XI42/XI581/MM6_g
+ N_XI42/XI581/NET21_XI42/XI581/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI613/MM6 N_NET305_XI42/XI613/MM6_d N_XI42/NET803_XI42/XI613/MM6_g
+ N_XI42/XI613/NET21_XI42/XI613/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI549/MM6 N_NET306_XI42/XI549/MM6_d N_XI42/NET245_XI42/XI549/MM6_g
+ N_XI42/XI549/NET21_XI42/XI549/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI629/MM6 N_NET307_XI42/XI629/MM6_d N_XI42/NET802_XI42/XI629/MM6_g
+ N_XI42/XI629/NET21_XI42/XI629/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI565/MM6 N_NET308_XI42/XI565/MM6_d N_XI42/NET375_XI42/XI565/MM6_g
+ N_XI42/XI565/NET21_XI42/XI565/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI597/MM6 N_NET309_XI42/XI597/MM6_d N_XI42/NET535_XI42/XI597/MM6_g
+ N_XI42/XI597/NET21_XI42/XI597/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI533/MM6 N_NET310_XI42/XI533/MM6_d N_XI42/NET180_XI42/XI533/MM6_g
+ N_XI42/XI533/NET21_XI42/XI533/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI644/MM6 N_NET311_XI42/XI644/MM6_d N_XI42/NET801_XI42/XI644/MM6_g
+ N_XI42/XI644/NET21_XI42/XI644/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI580/MM6 N_NET312_XI42/XI580/MM6_d N_XI42/NET455_XI42/XI580/MM6_g
+ N_XI42/XI580/NET21_XI42/XI580/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI612/MM6 N_NET313_XI42/XI612/MM6_d N_XI42/NET803_XI42/XI612/MM6_g
+ N_XI42/XI612/NET21_XI42/XI612/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI548/MM6 N_NET314_XI42/XI548/MM6_d N_XI42/NET245_XI42/XI548/MM6_g
+ N_XI42/XI548/NET21_XI42/XI548/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI628/MM6 N_NET315_XI42/XI628/MM6_d N_XI42/NET802_XI42/XI628/MM6_g
+ N_XI42/XI628/NET21_XI42/XI628/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI564/MM6 N_NET316_XI42/XI564/MM6_d N_XI42/NET375_XI42/XI564/MM6_g
+ N_XI42/XI564/NET21_XI42/XI564/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI596/MM6 N_NET317_XI42/XI596/MM6_d N_XI42/NET535_XI42/XI596/MM6_g
+ N_XI42/XI596/NET21_XI42/XI596/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI532/MM6 N_NET318_XI42/XI532/MM6_d N_XI42/NET180_XI42/XI532/MM6_g
+ N_XI42/XI532/NET21_XI42/XI532/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI643/MM6 N_NET319_XI42/XI643/MM6_d N_XI42/NET801_XI42/XI643/MM6_g
+ N_XI42/XI643/NET21_XI42/XI643/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI579/MM6 N_NET320_XI42/XI579/MM6_d N_XI42/NET455_XI42/XI579/MM6_g
+ N_XI42/XI579/NET21_XI42/XI579/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI611/MM6 N_NET321_XI42/XI611/MM6_d N_XI42/NET803_XI42/XI611/MM6_g
+ N_XI42/XI611/NET21_XI42/XI611/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI547/MM6 N_NET192_XI42/XI547/MM6_d N_XI42/NET245_XI42/XI547/MM6_g
+ N_XI42/XI547/NET21_XI42/XI547/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI627/MM6 N_NET193_XI42/XI627/MM6_d N_XI42/NET802_XI42/XI627/MM6_g
+ N_XI42/XI627/NET21_XI42/XI627/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI563/MM6 N_NET194_XI42/XI563/MM6_d N_XI42/NET375_XI42/XI563/MM6_g
+ N_XI42/XI563/NET21_XI42/XI563/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI595/MM6 N_NET195_XI42/XI595/MM6_d N_XI42/NET535_XI42/XI595/MM6_g
+ N_XI42/XI595/NET21_XI42/XI595/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI531/MM6 N_NET196_XI42/XI531/MM6_d N_XI42/NET180_XI42/XI531/MM6_g
+ N_XI42/XI531/NET21_XI42/XI531/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI642/MM6 N_NET197_XI42/XI642/MM6_d N_XI42/NET801_XI42/XI642/MM6_g
+ N_XI42/XI642/NET21_XI42/XI642/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI578/MM6 N_NET198_XI42/XI578/MM6_d N_XI42/NET455_XI42/XI578/MM6_g
+ N_XI42/XI578/NET21_XI42/XI578/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI610/MM6 N_NET199_XI42/XI610/MM6_d N_XI42/NET803_XI42/XI610/MM6_g
+ N_XI42/XI610/NET21_XI42/XI610/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI546/MM6 N_NET200_XI42/XI546/MM6_d N_XI42/NET245_XI42/XI546/MM6_g
+ N_XI42/XI546/NET21_XI42/XI546/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI626/MM6 N_NET331_XI42/XI626/MM6_d N_XI42/NET802_XI42/XI626/MM6_g
+ N_XI42/XI626/NET21_XI42/XI626/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI562/MM6 N_NET332_XI42/XI562/MM6_d N_XI42/NET375_XI42/XI562/MM6_g
+ N_XI42/XI562/NET21_XI42/XI562/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI594/MM6 N_NET203_XI42/XI594/MM6_d N_XI42/NET535_XI42/XI594/MM6_g
+ N_XI42/XI594/NET21_XI42/XI594/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI530/MM6 N_NET204_XI42/XI530/MM6_d N_XI42/NET180_XI42/XI530/MM6_g
+ N_XI42/XI530/NET21_XI42/XI530/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI641/MM6 N_NET205_XI42/XI641/MM6_d N_XI42/NET801_XI42/XI641/MM6_g
+ N_XI42/XI641/NET21_XI42/XI641/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI577/MM6 N_NET206_XI42/XI577/MM6_d N_XI42/NET455_XI42/XI577/MM6_g
+ N_XI42/XI577/NET21_XI42/XI577/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI609/MM6 N_NET207_XI42/XI609/MM6_d N_XI42/NET803_XI42/XI609/MM6_g
+ N_XI42/XI609/NET21_XI42/XI609/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI545/MM6 N_NET338_XI42/XI545/MM6_d N_XI42/NET245_XI42/XI545/MM6_g
+ N_XI42/XI545/NET21_XI42/XI545/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI625/MM6 N_NET339_XI42/XI625/MM6_d N_XI42/NET802_XI42/XI625/MM6_g
+ N_XI42/XI625/NET21_XI42/XI625/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI561/MM6 N_NET340_XI42/XI561/MM6_d N_XI42/NET375_XI42/XI561/MM6_g
+ N_XI42/XI561/NET21_XI42/XI561/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI593/MM6 N_NET211_XI42/XI593/MM6_d N_XI42/NET535_XI42/XI593/MM6_g
+ N_XI42/XI593/NET21_XI42/XI593/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI529/MM6 N_NET212_XI42/XI529/MM6_d N_XI42/NET180_XI42/XI529/MM6_g
+ N_XI42/XI529/NET21_XI42/XI529/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI640/MM6 N_NET214_XI42/XI640/MM6_d N_XI42/NET801_XI42/XI640/MM6_g
+ N_XI42/XI640/NET21_XI42/XI640/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI576/MM6 N_NET215_XI42/XI576/MM6_d N_XI42/NET455_XI42/XI576/MM6_g
+ N_XI42/XI576/NET21_XI42/XI576/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI608/MM6 N_NET216_XI42/XI608/MM6_d N_XI42/NET803_XI42/XI608/MM6_g
+ N_XI42/XI608/NET21_XI42/XI608/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI544/MM6 N_NET346_XI42/XI544/MM6_d N_XI42/NET245_XI42/XI544/MM6_g
+ N_XI42/XI544/NET21_XI42/XI544/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI624/MM6 N_NET347_XI42/XI624/MM6_d N_XI42/NET802_XI42/XI624/MM6_g
+ N_XI42/XI624/NET21_XI42/XI624/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI560/MM6 N_NET348_XI42/XI560/MM6_d N_XI42/NET375_XI42/XI560/MM6_g
+ N_XI42/XI560/NET21_XI42/XI560/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI592/MM6 N_NET349_XI42/XI592/MM6_d N_XI42/NET535_XI42/XI592/MM6_g
+ N_XI42/XI592/NET21_XI42/XI592/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI528/MM6 N_NET350_XI42/XI528/MM6_d N_XI42/NET180_XI42/XI528/MM6_g
+ N_XI42/XI528/NET21_XI42/XI528/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI639/MM6 N_NET351_XI42/XI639/MM6_d N_XI42/NET801_XI42/XI639/MM6_g
+ N_XI42/XI639/NET21_XI42/XI639/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI575/MM6 N_NET352_XI42/XI575/MM6_d N_XI42/NET455_XI42/XI575/MM6_g
+ N_XI42/XI575/NET21_XI42/XI575/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI607/MM6 N_NET224_XI42/XI607/MM6_d N_XI42/NET803_XI42/XI607/MM6_g
+ N_XI42/XI607/NET21_XI42/XI607/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI543/MM6 N_NET225_XI42/XI543/MM6_d N_XI42/NET245_XI42/XI543/MM6_g
+ N_XI42/XI543/NET21_XI42/XI543/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI623/MM6 N_NET226_XI42/XI623/MM6_d N_XI42/NET802_XI42/XI623/MM6_g
+ N_XI42/XI623/NET21_XI42/XI623/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI559/MM6 N_NET356_XI42/XI559/MM6_d N_XI42/NET375_XI42/XI559/MM6_g
+ N_XI42/XI559/NET21_XI42/XI559/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI591/MM6 N_NET357_XI42/XI591/MM6_d N_XI42/NET535_XI42/XI591/MM6_g
+ N_XI42/XI591/NET21_XI42/XI591/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI527/MM6 N_NET358_XI42/XI527/MM6_d N_XI42/NET180_XI42/XI527/MM6_g
+ N_XI42/XI527/NET21_XI42/XI527/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI638/MM6 N_NET230_XI42/XI638/MM6_d N_XI42/NET801_XI42/XI638/MM6_g
+ N_XI42/XI638/NET21_XI42/XI638/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI574/MM6 N_NET360_XI42/XI574/MM6_d N_XI42/NET455_XI42/XI574/MM6_g
+ N_XI42/XI574/NET21_XI42/XI574/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI606/MM6 N_NET361_XI42/XI606/MM6_d N_XI42/NET803_XI42/XI606/MM6_g
+ N_XI42/XI606/NET21_XI42/XI606/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI542/MM6 N_NET233_XI42/XI542/MM6_d N_XI42/NET245_XI42/XI542/MM6_g
+ N_XI42/XI542/NET21_XI42/XI542/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI622/MM6 N_NET234_XI42/XI622/MM6_d N_XI42/NET802_XI42/XI622/MM6_g
+ N_XI42/XI622/NET21_XI42/XI622/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI558/MM6 N_NET235_XI42/XI558/MM6_d N_XI42/NET375_XI42/XI558/MM6_g
+ N_XI42/XI558/NET21_XI42/XI558/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI590/MM6 N_NET365_XI42/XI590/MM6_d N_XI42/NET535_XI42/XI590/MM6_g
+ N_XI42/XI590/NET21_XI42/XI590/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI526/MM6 N_NET366_XI42/XI526/MM6_d N_XI42/NET180_XI42/XI526/MM6_g
+ N_XI42/XI526/NET21_XI42/XI526/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI637/MM6 N_NET367_XI42/XI637/MM6_d N_XI42/NET801_XI42/XI637/MM6_g
+ N_XI42/XI637/NET21_XI42/XI637/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI573/MM6 N_NET368_XI42/XI573/MM6_d N_XI42/NET455_XI42/XI573/MM6_g
+ N_XI42/XI573/NET21_XI42/XI573/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI605/MM6 N_NET369_XI42/XI605/MM6_d N_XI42/NET803_XI42/XI605/MM6_g
+ N_XI42/XI605/NET21_XI42/XI605/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI541/MM6 N_NET370_XI42/XI541/MM6_d N_XI42/NET245_XI42/XI541/MM6_g
+ N_XI42/XI541/NET21_XI42/XI541/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI621/MM6 N_NET371_XI42/XI621/MM6_d N_XI42/NET802_XI42/XI621/MM6_g
+ N_XI42/XI621/NET21_XI42/XI621/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI557/MM6 N_NET242_XI42/XI557/MM6_d N_XI42/NET375_XI42/XI557/MM6_g
+ N_XI42/XI557/NET21_XI42/XI557/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI589/MM6 N_NET373_XI42/XI589/MM6_d N_XI42/NET535_XI42/XI589/MM6_g
+ N_XI42/XI589/NET21_XI42/XI589/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI525/MM6 N_NET244_XI42/XI525/MM6_d N_XI42/NET180_XI42/XI525/MM6_g
+ N_XI42/XI525/NET21_XI42/XI525/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI636/MM6 N_NET375_XI42/XI636/MM6_d N_XI42/NET801_XI42/XI636/MM6_g
+ N_XI42/XI636/NET21_XI42/XI636/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI572/MM6 N_NET376_XI42/XI572/MM6_d N_XI42/NET455_XI42/XI572/MM6_g
+ N_XI42/XI572/NET21_XI42/XI572/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI604/MM6 N_NET377_XI42/XI604/MM6_d N_XI42/NET803_XI42/XI604/MM6_g
+ N_XI42/XI604/NET21_XI42/XI604/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI540/MM6 N_NET378_XI42/XI540/MM6_d N_XI42/NET245_XI42/XI540/MM6_g
+ N_XI42/XI540/NET21_XI42/XI540/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI620/MM6 N_NET379_XI42/XI620/MM6_d N_XI42/NET802_XI42/XI620/MM6_g
+ N_XI42/XI620/NET21_XI42/XI620/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI556/MM6 N_NET380_XI42/XI556/MM6_d N_XI42/NET375_XI42/XI556/MM6_g
+ N_XI42/XI556/NET21_XI42/XI556/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI588/MM6 N_NET381_XI42/XI588/MM6_d N_XI42/NET535_XI42/XI588/MM6_g
+ N_XI42/XI588/NET21_XI42/XI588/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI524/MM6 N_NET382_XI42/XI524/MM6_d N_XI42/NET180_XI42/XI524/MM6_g
+ N_XI42/XI524/NET21_XI42/XI524/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI635/MM6 N_NET383_XI42/XI635/MM6_d N_XI42/NET801_XI42/XI635/MM6_g
+ N_XI42/XI635/NET21_XI42/XI635/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI571/MM6 N_NET384_XI42/XI571/MM6_d N_XI42/NET455_XI42/XI571/MM6_g
+ N_XI42/XI571/NET21_XI42/XI571/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI603/MM6 N_NET385_XI42/XI603/MM6_d N_XI42/NET803_XI42/XI603/MM6_g
+ N_XI42/XI603/NET21_XI42/XI603/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI539/MM6 N_NET256_XI42/XI539/MM6_d N_XI42/NET245_XI42/XI539/MM6_g
+ N_XI42/XI539/NET21_XI42/XI539/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI619/MM6 N_NET387_XI42/XI619/MM6_d N_XI42/NET802_XI42/XI619/MM6_g
+ N_XI42/XI619/NET21_XI42/XI619/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI555/MM6 N_NET388_XI42/XI555/MM6_d N_XI42/NET375_XI42/XI555/MM6_g
+ N_XI42/XI555/NET21_XI42/XI555/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI587/MM6 N_NET389_XI42/XI587/MM6_d N_XI42/NET535_XI42/XI587/MM6_g
+ N_XI42/XI587/NET21_XI42/XI587/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI523/MM6 N_NET390_XI42/XI523/MM6_d N_XI42/NET180_XI42/XI523/MM6_g
+ N_XI42/XI523/NET21_XI42/XI523/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI634/MM6 N_NET391_XI42/XI634/MM6_d N_XI42/NET801_XI42/XI634/MM6_g
+ N_XI42/XI634/NET21_XI42/XI634/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI570/MM6 N_NET262_XI42/XI570/MM6_d N_XI42/NET455_XI42/XI570/MM6_g
+ N_XI42/XI570/NET21_XI42/XI570/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI602/MM6 N_NET263_XI42/XI602/MM6_d N_XI42/NET803_XI42/XI602/MM6_g
+ N_XI42/XI602/NET21_XI42/XI602/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI538/MM6 N_NET264_XI42/XI538/MM6_d N_XI42/NET245_XI42/XI538/MM6_g
+ N_XI42/XI538/NET21_XI42/XI538/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI618/MM6 N_NET265_XI42/XI618/MM6_d N_XI42/NET802_XI42/XI618/MM6_g
+ N_XI42/XI618/NET21_XI42/XI618/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI554/MM6 N_NET396_XI42/XI554/MM6_d N_XI42/NET375_XI42/XI554/MM6_g
+ N_XI42/XI554/NET21_XI42/XI554/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI586/MM6 N_NET267_XI42/XI586/MM6_d N_XI42/NET535_XI42/XI586/MM6_g
+ N_XI42/XI586/NET21_XI42/XI586/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI522/MM6 N_NET268_XI42/XI522/MM6_d N_XI42/NET180_XI42/XI522/MM6_g
+ N_XI42/XI522/NET21_XI42/XI522/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI633/MM6 N_NET269_XI42/XI633/MM6_d N_XI42/NET801_XI42/XI633/MM6_g
+ N_XI42/XI633/NET21_XI42/XI633/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI569/MM6 N_NET270_XI42/XI569/MM6_d N_XI42/NET455_XI42/XI569/MM6_g
+ N_XI42/XI569/NET21_XI42/XI569/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI601/MM6 N_NET401_XI42/XI601/MM6_d N_XI42/NET803_XI42/XI601/MM6_g
+ N_XI42/XI601/NET21_XI42/XI601/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI537/MM6 N_NET272_XI42/XI537/MM6_d N_XI42/NET245_XI42/XI537/MM6_g
+ N_XI42/XI537/NET21_XI42/XI537/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI617/MM6 N_NET273_XI42/XI617/MM6_d N_XI42/NET802_XI42/XI617/MM6_g
+ N_XI42/XI617/NET21_XI42/XI617/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI553/MM6 N_NET404_XI42/XI553/MM6_d N_XI42/NET375_XI42/XI553/MM6_g
+ N_XI42/XI553/NET21_XI42/XI553/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI585/MM6 N_NET405_XI42/XI585/MM6_d N_XI42/NET535_XI42/XI585/MM6_g
+ N_XI42/XI585/NET21_XI42/XI585/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI42/XI521/MM6 N_XI42/NET0388_XI42/XI521/MM6_d N_XI42/NET180_XI42/XI521/MM6_g
+ N_XI42/XI521/NET21_XI42/XI521/MM6_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07
+ W=4.7e-07 AD=2.397e-13 AS=7.05e-14 PD=1.49e-06 PS=3e-07
mXI39/MM16 N_NET0380_XI39/MM16_d N_NET070_XI39/MM16_g N_VDD_XI39/MM16_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI29/XI0/MM31 N_NET064_XI29/XI0/MM31_d N_NET470_XI29/XI0/MM31_g
+ N_NET0380_XI29/XI0/MM31_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI29/XI0/XI8/MM0 N_XI29/XI0/NET195_XI29/XI0/XI8/MM0_d
+ N_NET470_XI29/XI0/XI8/MM0_g N_VDD_XI29/XI0/XI8/MM0_s N_VDD_XI29/XI0/XI8/MM0_b
+ P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI29/XI0/MM32 N_NET064_XI29/XI0/MM32_d N_NET469_XI29/XI0/MM32_g
+ N_NET474_XI29/XI0/MM32_s N_VDD_XI29/XI0/MM32_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI29/XI0/XI9/MM0 N_XI29/XI0/NET199_XI29/XI0/XI9/MM0_d
+ N_NET469_XI29/XI0/XI9/MM0_g N_VDD_XI29/XI0/XI9/MM0_s N_VDD_XI29/XI0/XI9/MM0_b
+ P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI39/MM17 N_NET474_XI39/MM17_d N_NET070_XI39/MM17_g N_VDD_XI39/MM17_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI29/XI0/MM33 N_NET064_XI29/XI0/MM33_d N_NET468_XI29/XI0/MM33_g
+ N_NET475_XI29/XI0/MM33_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI29/XI0/XI10/MM0 N_XI29/XI0/NET223_XI29/XI0/XI10/MM0_d
+ N_NET468_XI29/XI0/XI10/MM0_g N_VDD_XI29/XI0/XI10/MM0_s
+ N_VDD_XI29/XI0/XI8/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=2.303e-13
+ PD=1.45e-06 PS=1.45e-06
mXI29/XI0/MM34 N_NET064_XI29/XI0/MM34_d N_NET467_XI29/XI0/MM34_g
+ N_NET476_XI29/XI0/MM34_s N_VDD_XI29/XI0/MM32_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI29/XI0/XI11/MM0 N_XI29/XI0/NET215_XI29/XI0/XI11/MM0_d
+ N_NET467_XI29/XI0/XI11/MM0_g N_VDD_XI29/XI0/XI11/MM0_s
+ N_VDD_XI29/XI0/XI9/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=2.303e-13
+ PD=1.45e-06 PS=1.45e-06
mXI39/MM18 N_NET475_XI39/MM18_d N_NET070_XI39/MM18_g N_VDD_XI39/MM18_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI39/MM19 N_NET476_XI39/MM19_d N_NET070_XI39/MM19_g N_VDD_XI39/MM19_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI57/XI1/MM3 N_XI57/NET12_XI57/XI1/MM3_d N_NET068_XI57/XI1/MM3_g
+ N_VDD_XI57/XI1/MM3_s N_VDD_XI57/XI1/MM3_b P_18 L=1.8e-07 W=4.7e-07 AD=2.35e-13
+ AS=1.7625e-13 PD=1.47e-06 PS=7.5e-07
mXI57/XI1/MM2 N_XI57/NET12_XI57/XI1/MM2_d N_NET061_XI57/XI1/MM2_g
+ N_VDD_XI57/XI1/MM2_s N_VDD_XI57/XI1/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.3735e-13 AS=1.7625e-13 PD=1.48e-06 PS=7.5e-07
mXI57/XI1/MM1 N_NET061_XI57/XI1/MM1_d N_XI57/NET12_XI57/XI1/MM1_g
+ N_VDD_XI57/XI1/MM1_s N_VDD_XI57/XI1/MM3_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.3735e-13 AS=1.7625e-13 PD=1.48e-06 PS=7.5e-07
mXI57/XI1/MM0 N_NET061_XI57/XI1/MM0_d N_NET068_XI57/XI1/MM0_g
+ N_VDD_XI57/XI1/MM0_s N_VDD_XI57/XI1/MM3_b P_18 L=1.8e-07 W=4.7e-07 AD=2.35e-13
+ AS=1.7625e-13 PD=1.47e-06 PS=7.5e-07
mXI39/MM20 N_NET414_XI39/MM20_d N_NET070_XI39/MM20_g N_VDD_XI39/MM20_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI29/XI0/MM35 N_NET064_XI29/XI0/MM35_d N_NET466_XI29/XI0/MM35_g
+ N_NET414_XI29/XI0/MM35_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI29/XI0/XI12/MM0 N_XI29/XI0/NET211_XI29/XI0/XI12/MM0_d
+ N_NET466_XI29/XI0/XI12/MM0_g N_VDD_XI29/XI0/XI12/MM0_s
+ N_VDD_XI29/XI0/XI8/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=2.303e-13
+ PD=1.45e-06 PS=1.45e-06
mXI29/XI0/MM36 N_NET064_XI29/XI0/MM36_d N_NET465_XI29/XI0/MM36_g
+ N_NET415_XI29/XI0/MM36_s N_VDD_XI29/XI0/MM32_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI29/XI0/XI13/MM0 N_XI29/XI0/NET203_XI29/XI0/XI13/MM0_d
+ N_NET465_XI29/XI0/XI13/MM0_g N_VDD_XI29/XI0/XI13/MM0_s
+ N_VDD_XI29/XI0/XI9/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=2.303e-13
+ PD=1.45e-06 PS=1.45e-06
mXI39/MM21 N_NET415_XI39/MM21_d N_NET070_XI39/MM21_g N_VDD_XI39/MM21_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI29/XI0/MM37 N_NET064_XI29/XI0/MM37_d N_NET464_XI29/XI0/MM37_g
+ N_NET416_XI29/XI0/MM37_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI29/XI0/XI14/MM0 N_XI29/XI0/NET219_XI29/XI0/XI14/MM0_d
+ N_NET464_XI29/XI0/XI14/MM0_g N_VDD_XI29/XI0/XI14/MM0_s
+ N_VDD_XI29/XI0/XI8/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=2.303e-13
+ PD=1.45e-06 PS=1.45e-06
mXI29/XI0/MM38 N_NET064_XI29/XI0/MM38_d N_NET463_XI29/XI0/MM38_g
+ N_NET417_XI29/XI0/MM38_s N_VDD_XI29/XI0/MM32_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI29/XI0/XI15/MM0 N_XI29/XI0/NET207_XI29/XI0/XI15/MM0_d
+ N_NET463_XI29/XI0/XI15/MM0_g N_VDD_XI29/XI0/XI15/MM0_s
+ N_VDD_XI29/XI0/XI9/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=2.303e-13
+ PD=1.45e-06 PS=1.45e-06
mXI39/MM22 N_NET416_XI39/MM22_d N_NET070_XI39/MM22_g N_VDD_XI39/MM22_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI54/XI1/XI6/MM0 N_XI54/XI1/NET2_XI54/XI1/XI6/MM0_d N_NET061_XI54/XI1/XI6/MM0_g
+ N_VDD_XI54/XI1/XI6/MM0_s N_VDD_XI57/XI1/MM3_b P_18 L=1.8e-07 W=1.85e-06
+ AD=9.435e-13 AS=9.435e-13 PD=2.87e-06 PS=2.87e-06
mXI39/MM23 N_NET417_XI39/MM23_d N_NET070_XI39/MM23_g N_VDD_XI39/MM23_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI29/XI1/MM31 N_NET065_XI29/XI1/MM31_d N_NET470_XI29/XI1/MM31_g
+ N_NET481_XI29/XI1/MM31_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI29/XI1/XI8/MM0 N_XI29/XI1/NET195_XI29/XI1/XI8/MM0_d
+ N_NET470_XI29/XI1/XI8/MM0_g N_VDD_XI29/XI1/XI8/MM0_s N_VDD_XI29/XI0/XI8/MM0_b
+ P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI29/XI1/MM32 N_NET065_XI29/XI1/MM32_d N_NET469_XI29/XI1/MM32_g
+ N_NET482_XI29/XI1/MM32_s N_VDD_XI29/XI0/MM32_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI29/XI1/XI9/MM0 N_XI29/XI1/NET199_XI29/XI1/XI9/MM0_d
+ N_NET469_XI29/XI1/XI9/MM0_g N_VDD_XI29/XI1/XI9/MM0_s N_VDD_XI29/XI0/XI9/MM0_b
+ P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI39/MM24 N_NET481_XI39/MM24_d N_NET070_XI39/MM24_g N_VDD_XI39/MM24_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI54/XI1/XI8/XI3/MM1 N_XI54/XI1/XI8/NET12_XI54/XI1/XI8/XI3/MM1_d
+ N_XI54/XI1/NET2_XI54/XI1/XI8/XI3/MM1_g N_VDD_XI54/XI1/XI8/XI3/MM1_s
+ N_VDD_XI57/XI1/MM3_b P_18 L=1.8e-07 W=4.7e-07 AD=1.68025e-13 AS=2.303e-13
+ PD=7.15e-07 PS=1.45e-06
mXI54/XI1/XI7/XI3/MM1 N_XI54/XI1/XI7/NET12_XI54/XI1/XI7/XI3/MM1_d
+ N_NET061_XI54/XI1/XI7/XI3/MM1_g N_VDD_XI54/XI1/XI7/XI3/MM1_s
+ N_VDD_XI54/XI1/XI7/XI3/MM1_b P_18 L=1.8e-07 W=4.7e-07 AD=1.68025e-13
+ AS=2.5145e-13 PD=7.15e-07 PS=1.54e-06
mXI39/MM25 N_NET482_XI39/MM25_d N_NET070_XI39/MM25_g N_VDD_XI39/MM25_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI54/XI1/XI8/XI3/MM0 N_XI54/XI1/XI8/NET12_XI54/XI1/XI8/XI3/MM0_d
+ N_NET068_XI54/XI1/XI8/XI3/MM0_g N_VDD_XI54/XI1/XI8/XI3/MM0_s
+ N_VDD_XI57/XI1/MM3_b P_18 L=1.8e-07 W=4.7e-07 AD=1.68025e-13 AS=2.3265e-13
+ PD=7.15e-07 PS=1.46e-06
mXI54/XI1/XI7/XI3/MM0 N_XI54/XI1/XI7/NET12_XI54/XI1/XI7/XI3/MM0_d
+ N_NET068_XI54/XI1/XI7/XI3/MM0_g N_VDD_XI54/XI1/XI7/XI3/MM0_s
+ N_VDD_XI54/XI1/XI7/XI3/MM1_b P_18 L=1.8e-07 W=4.7e-07 AD=1.68025e-13
+ AS=2.3265e-13 PD=7.15e-07 PS=1.46e-06
mXI29/XI1/MM33 N_NET065_XI29/XI1/MM33_d N_NET468_XI29/XI1/MM33_g
+ N_NET420_XI29/XI1/MM33_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI29/XI1/XI10/MM0 N_XI29/XI1/NET223_XI29/XI1/XI10/MM0_d
+ N_NET468_XI29/XI1/XI10/MM0_g N_VDD_XI29/XI1/XI10/MM0_s
+ N_VDD_XI29/XI0/XI8/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=2.303e-13
+ PD=1.45e-06 PS=1.45e-06
mXI29/XI1/MM34 N_NET065_XI29/XI1/MM34_d N_NET467_XI29/XI1/MM34_g
+ N_NET421_XI29/XI1/MM34_s N_VDD_XI29/XI0/MM32_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI29/XI1/XI11/MM0 N_XI29/XI1/NET215_XI29/XI1/XI11/MM0_d
+ N_NET467_XI29/XI1/XI11/MM0_g N_VDD_XI29/XI1/XI11/MM0_s
+ N_VDD_XI29/XI0/XI9/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=2.303e-13
+ PD=1.45e-06 PS=1.45e-06
mXI39/MM26 N_NET420_XI39/MM26_d N_NET070_XI39/MM26_g N_VDD_XI39/MM26_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI39/MM27 N_NET421_XI39/MM27_d N_NET070_XI39/MM27_g N_VDD_XI39/MM27_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI54/XI1/XI8/XI2/MM0 N_XI54/XI1/NET9_XI54/XI1/XI8/XI2/MM0_d
+ N_XI54/XI1/XI8/NET12_XI54/XI1/XI8/XI2/MM0_g N_VDD_XI54/XI1/XI8/XI2/MM0_s
+ N_VDD_XI57/XI1/MM3_b P_18 L=1.8e-07 W=1.85e-06 AD=9.435e-13 AS=9.435e-13
+ PD=2.87e-06 PS=2.87e-06
mXI54/XI1/XI7/XI2/MM0 N_XI54/XI1/NET10_XI54/XI1/XI7/XI2/MM0_d
+ N_XI54/XI1/XI7/NET12_XI54/XI1/XI7/XI2/MM0_g N_VDD_XI54/XI1/XI7/XI2/MM0_s
+ N_VDD_XI54/XI1/XI7/XI3/MM1_b P_18 L=1.8e-07 W=1.85e-06 AD=9.435e-13
+ AS=9.435e-13 PD=2.87e-06 PS=2.87e-06
mXI29/XI1/MM35 N_NET065_XI29/XI1/MM35_d N_NET466_XI29/XI1/MM35_g
+ N_NET485_XI29/XI1/MM35_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI29/XI1/XI12/MM0 N_XI29/XI1/NET211_XI29/XI1/XI12/MM0_d
+ N_NET466_XI29/XI1/XI12/MM0_g N_VDD_XI29/XI1/XI12/MM0_s
+ N_VDD_XI29/XI0/XI8/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=2.303e-13
+ PD=1.45e-06 PS=1.45e-06
mXI29/XI1/MM36 N_NET065_XI29/XI1/MM36_d N_NET465_XI29/XI1/MM36_g
+ N_NET486_XI29/XI1/MM36_s N_VDD_XI29/XI0/MM32_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI29/XI1/XI13/MM0 N_XI29/XI1/NET203_XI29/XI1/XI13/MM0_d
+ N_NET465_XI29/XI1/XI13/MM0_g N_VDD_XI29/XI1/XI13/MM0_s
+ N_VDD_XI29/XI0/XI9/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=2.303e-13
+ PD=1.45e-06 PS=1.45e-06
mXI39/MM28 N_NET485_XI39/MM28_d N_NET070_XI39/MM28_g N_VDD_XI39/MM28_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI39/MM29 N_NET486_XI39/MM29_d N_NET070_XI39/MM29_g N_VDD_XI39/MM29_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI54/XI1/XI10/MM6 N_XI54/XI1/XI10/NET21_XI54/XI1/XI10/MM6_d
+ N_XI54/XI1/NET9_XI54/XI1/XI10/MM6_g N_VDD_XI54/XI1/XI10/MM6_s
+ N_VDD_XI57/XI1/MM3_b P_18 L=1.8e-07 W=4.7e-07 AD=1.68025e-13 AS=2.303e-13
+ PD=7.15e-07 PS=1.45e-06
mXI54/XI1/XI9/MM6 N_XI54/XI1/XI9/NET21_XI54/XI1/XI9/MM6_d
+ N_DOUT<1>_XI54/XI1/XI9/MM6_g N_VDD_XI54/XI1/XI9/MM6_s
+ N_VDD_XI54/XI1/XI7/XI3/MM1_b P_18 L=1.8e-07 W=4.7e-07 AD=1.68025e-13
+ AS=2.5145e-13 PD=7.15e-07 PS=1.54e-06
mXI54/XI1/XI10/MM7 N_DOUT<1>_XI54/XI1/XI10/MM7_d
+ N_XI54/NET16_XI54/XI1/XI10/MM7_g N_XI54/XI1/XI10/NET21_XI54/XI1/XI10/MM7_s
+ N_VDD_XI57/XI1/MM3_b P_18 L=1.8e-07 W=4.7e-07 AD=2.3265e-13 AS=1.68025e-13
+ PD=1.46e-06 PS=7.15e-07
mXI54/XI1/XI9/MM7 N_XI54/NET16_XI54/XI1/XI9/MM7_d
+ N_XI54/XI1/NET10_XI54/XI1/XI9/MM7_g N_XI54/XI1/XI9/NET21_XI54/XI1/XI9/MM7_s
+ N_VDD_XI54/XI1/XI7/XI3/MM1_b P_18 L=1.8e-07 W=4.7e-07 AD=2.3265e-13
+ AS=1.68025e-13 PD=1.46e-06 PS=7.15e-07
mXI29/XI1/MM37 N_NET065_XI29/XI1/MM37_d N_NET464_XI29/XI1/MM37_g
+ N_NET487_XI29/XI1/MM37_s N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI29/XI1/XI14/MM0 N_XI29/XI1/NET219_XI29/XI1/XI14/MM0_d
+ N_NET464_XI29/XI1/XI14/MM0_g N_VDD_XI29/XI1/XI14/MM0_s
+ N_VDD_XI29/XI0/XI8/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=2.303e-13
+ PD=1.45e-06 PS=1.45e-06
mXI29/XI1/MM38 N_NET065_XI29/XI1/MM38_d N_NET463_XI29/XI1/MM38_g
+ N_NET0395_XI29/XI1/MM38_s N_VDD_XI29/XI0/MM32_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI29/XI1/XI15/MM0 N_XI29/XI1/NET207_XI29/XI1/XI15/MM0_d
+ N_NET463_XI29/XI1/XI15/MM0_g N_VDD_XI29/XI1/XI15/MM0_s
+ N_VDD_XI29/XI0/XI9/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=2.303e-13
+ PD=1.45e-06 PS=1.45e-06
mXI39/MM30 N_NET487_XI39/MM30_d N_NET070_XI39/MM30_g N_VDD_XI39/MM30_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXI39/MM31 N_NET0395_XI39/MM31_d N_NET070_XI39/MM31_g N_VDD_XI39/MM31_s
+ N_VDD_XI42/XI649/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
c_1 XI39/NET5650 0 0.15106f
c_2 XI39/NET5466 0 0.150863f
c_3 XI39/NET5718 0 0.150863f
c_4 XI39/NET3574 0 0.150863f
c_5 XI39/NET5210 0 0.150863f
c_6 XI39/NET5398 0 0.150863f
c_7 XI39/NET5142 0 0.150863f
c_8 XI39/NET4954 0 0.150863f
c_9 XI39/NET3930 0 0.150863f
c_10 XI39/NET4118 0 0.150863f
c_11 XI39/NET3862 0 0.150863f
c_12 XI39/NET3674 0 0.150863f
c_13 XI39/NET4374 0 0.150863f
c_14 XI39/NET4186 0 0.150863f
c_15 XI39/NET4442 0 0.150863f
c_16 XI39/NET4630 0 0.150863f
c_17 XI39/NET6126 0 0.150863f
c_18 XI39/NET7462 0 0.150863f
c_19 XI39/NET6058 0 0.150863f
c_20 XI39/NET5870 0 0.150863f
c_21 XI39/NET7142 0 0.150863f
c_22 XI39/NET7530 0 0.150863f
c_23 XI39/NET7210 0 0.150863f
c_24 XI39/NET7022 0 0.150863f
c_25 XI39/NET6418 0 0.150863f
c_26 XI39/NET6230 0 0.150863f
c_27 XI39/NET6486 0 0.150863f
c_28 XI39/NET6674 0 0.150863f
c_29 XI39/NET4698 0 0.150863f
c_30 XI39/NET4886 0 0.150863f
c_31 XI39/NET6930 0 0.150863f
c_32 XI39/NET6770 0 0.150863f
c_33 XI39/NET8922 0 0.150863f
c_34 XI39/NET9106 0 0.150863f
c_35 XI39/NET8854 0 0.150863f
c_36 XI39/NET8666 0 0.150863f
c_37 XI39/NET9362 0 0.150863f
c_38 XI39/NET9174 0 0.150863f
c_39 XI39/NET9430 0 0.150863f
c_40 XI39/NET9618 0 0.150863f
c_41 XI39/NET8342 0 0.150863f
c_42 XI39/NET8154 0 0.150863f
c_43 XI39/NET8410 0 0.150863f
c_44 XI39/NET8598 0 0.150863f
c_45 XI39/NET7898 0 0.150863f
c_46 XI39/NET8086 0 0.150863f
c_47 XI39/NET7830 0 0.150863f
c_48 XI39/NET7642 0 0.150863f
c_49 XI39/NET10746 0 0.150863f
c_50 XI39/NET11206 0 0.150863f
c_51 XI39/NET10814 0 0.150863f
c_52 XI39/NET11002 0 0.150863f
c_53 XI39/NET11526 0 0.150863f
c_54 XI39/NET11138 0 0.150863f
c_55 XI39/NET11458 0 0.150863f
c_56 XI39/NET11646 0 0.150863f
c_57 XI39/NET10458 0 0.150863f
c_58 XI39/NET10638 0 0.150863f
c_59 XI39/NET10390 0 0.150863f
c_60 XI39/NET10210 0 0.150863f
c_61 XI39/NET9874 0 0.150863f
c_62 XI39/NET9694 0 0.150863f
c_63 XI39/NET9946 0 0.150863f
c_64 XI39/NET10098 0 0.149709f
c_65 XI39/NET5590 0 0.180473f
c_66 XI39/NET5530 0 0.176433f
c_67 XI39/NET5782 0 0.176433f
c_68 XI39/NET3542 0 0.176433f
c_69 XI39/NET5274 0 0.176433f
c_70 XI39/NET5334 0 0.176433f
c_71 XI39/NET5078 0 0.176433f
c_72 XI39/NET5018 0 0.176433f
c_73 XI39/NET3994 0 0.18066f
c_74 XI39/NET4054 0 0.176433f
c_75 XI39/NET3798 0 0.176433f
c_76 XI39/NET3738 0 0.176433f
c_77 XI39/NET4310 0 0.176433f
c_78 XI39/NET4250 0 0.176433f
c_79 XI39/NET4506 0 0.176433f
c_80 XI39/NET4566 0 0.176433f
c_81 XI39/NET7338 0 0.18066f
c_82 XI39/NET7398 0 0.176433f
c_83 XI39/NET5994 0 0.176433f
c_84 XI39/NET5934 0 0.176433f
c_85 XI39/NET7078 0 0.176433f
c_86 XI39/NET7578 0 0.176433f
c_87 XI39/NET7274 0 0.176433f
c_88 XI39/NET7310 0 0.176433f
c_89 XI39/NET6354 0 0.18066f
c_90 XI39/NET6294 0 0.176433f
c_91 XI39/NET6550 0 0.176433f
c_92 XI39/NET6610 0 0.176433f
c_93 XI39/NET4762 0 0.176433f
c_94 XI39/NET4822 0 0.176433f
c_95 XI39/NET6866 0 0.176433f
c_96 XI39/NET6802 0 0.176433f
c_97 XI39/NET8982 0 0.18066f
c_98 XI39/NET9042 0 0.176433f
c_99 XI39/NET8790 0 0.176433f
c_100 XI39/NET8730 0 0.176433f
c_101 XI39/NET9298 0 0.176433f
c_102 XI39/NET9238 0 0.176433f
c_103 XI39/NET9494 0 0.176433f
c_104 XI39/NET9554 0 0.176433f
c_105 XI39/NET8278 0 0.18066f
c_106 XI39/NET8218 0 0.176433f
c_107 XI39/NET8474 0 0.176433f
c_108 XI39/NET8534 0 0.176433f
c_109 XI39/NET7962 0 0.176433f
c_110 XI39/NET8022 0 0.176433f
c_111 XI39/NET7766 0 0.176433f
c_112 XI39/NET7706 0 0.176433f
c_113 XI39/NET11290 0 0.18066f
c_114 XI39/NET11270 0 0.176433f
c_115 XI39/NET10878 0 0.176433f
c_116 XI39/NET10938 0 0.176433f
c_117 XI39/NET11582 0 0.176433f
c_118 XI39/NET11074 0 0.176433f
c_119 XI39/NET11394 0 0.176433f
c_120 XI39/NET11670 0 0.176433f
c_121 XI39/NET10518 0 0.18066f
c_122 XI39/NET10578 0 0.176433f
c_123 XI39/NET10330 0 0.176433f
c_124 XI39/NET10270 0 0.176433f
c_125 XI39/NET9814 0 0.176433f
c_126 XI39/NET9754 0 0.176433f
c_127 XI39/NET10006 0 0.176433f
c_128 XI39/NET10130 0 0.176433f
c_129 XI39/NET5594 0 0.176433f
c_130 XI39/NET5410 0 0.176433f
c_131 XI39/NET5662 0 0.176433f
c_132 XI39/NET3566 0 0.176433f
c_133 XI39/NET5154 0 0.176433f
c_134 XI39/NET5342 0 0.176433f
c_135 XI39/NET5086 0 0.176433f
c_136 XI39/NET4898 0 0.176433f
c_137 XI39/NET3874 0 0.176433f
c_138 XI39/NET4062 0 0.176433f
c_139 XI39/NET3806 0 0.176433f
c_140 XI39/NET3618 0 0.176433f
c_141 XI39/NET4318 0 0.176433f
c_142 XI39/NET4130 0 0.176433f
c_143 XI39/NET4386 0 0.176433f
c_144 XI39/NET4574 0 0.176433f
c_145 XI39/NET6070 0 0.176433f
c_146 XI39/NET7406 0 0.176433f
c_147 XI39/NET6002 0 0.176433f
c_148 XI39/NET5814 0 0.176433f
c_149 XI39/NET7086 0 0.176433f
c_150 XI39/NET7474 0 0.176433f
c_151 XI39/NET7154 0 0.176433f
c_152 XI39/NET6966 0 0.176433f
c_153 XI39/NET6362 0 0.176433f
c_154 XI39/NET6174 0 0.176433f
c_155 XI39/NET6430 0 0.176433f
c_156 XI39/NET6618 0 0.176433f
c_157 XI39/NET4642 0 0.176433f
c_158 XI39/NET4830 0 0.176433f
c_159 XI39/NET6874 0 0.176433f
c_160 XI39/NET6714 0 0.176433f
c_161 XI39/NET8866 0 0.176433f
c_162 XI39/NET9050 0 0.176433f
c_163 XI39/NET8798 0 0.176433f
c_164 XI39/NET8610 0 0.176433f
c_165 XI39/NET9306 0 0.176433f
c_166 XI39/NET9118 0 0.176433f
c_167 XI39/NET9374 0 0.176433f
c_168 XI39/NET9562 0 0.176433f
c_169 XI39/NET8286 0 0.176433f
c_170 XI39/NET8098 0 0.176433f
c_171 XI39/NET8354 0 0.176433f
c_172 XI39/NET8542 0 0.176433f
c_173 XI39/NET7842 0 0.176433f
c_174 XI39/NET8030 0 0.176433f
c_175 XI39/NET7774 0 0.176433f
c_176 XI39/NET7586 0 0.176433f
c_177 XI39/NET10690 0 0.176433f
c_178 XI39/NET11150 0 0.176433f
c_179 XI39/NET10758 0 0.176433f
c_180 XI39/NET10946 0 0.176433f
c_181 XI39/NET11470 0 0.176433f
c_182 XI39/NET11082 0 0.176433f
c_183 XI39/NET11402 0 0.176433f
c_184 XI39/NET11590 0 0.176433f
c_185 XI39/NET10402 0 0.176433f
c_186 XI39/NET10582 0 0.176433f
c_187 XI39/NET10334 0 0.176433f
c_188 XI39/NET10154 0 0.176433f
c_189 XI39/NET9818 0 0.176433f
c_190 XI39/NET9638 0 0.176433f
c_191 XI39/NET9890 0 0.176433f
c_192 XI39/NET10066 0 0.176434f
c_193 XI39/NET5558 0 0.180473f
c_194 XI39/NET5482 0 0.176433f
c_195 XI39/NET5734 0 0.176433f
c_196 XI39/NET3494 0 0.176433f
c_197 XI39/NET5226 0 0.176433f
c_198 XI39/NET5286 0 0.176433f
c_199 XI39/NET5030 0 0.176433f
c_200 XI39/NET4970 0 0.176433f
c_201 XI39/NET3946 0 0.18066f
c_202 XI39/NET4006 0 0.176433f
c_203 XI39/NET3750 0 0.176433f
c_204 XI39/NET3690 0 0.176433f
c_205 XI39/NET4262 0 0.176433f
c_206 XI39/NET4202 0 0.176433f
c_207 XI39/NET4458 0 0.176433f
c_208 XI39/NET4518 0 0.176433f
c_209 XI39/NET6142 0 0.18066f
c_210 XI39/NET7350 0 0.176433f
c_211 XI39/NET5946 0 0.176433f
c_212 XI39/NET5886 0 0.176433f
c_213 XI39/NET7030 0 0.176433f
c_214 XI39/NET5798 0 0.176433f
c_215 XI39/NET7226 0 0.176433f
c_216 XI39/NET6950 0 0.176433f
c_217 XI39/NET6306 0 0.18066f
c_218 XI39/NET6246 0 0.176433f
c_219 XI39/NET6502 0 0.176433f
c_220 XI39/NET6562 0 0.176433f
c_221 XI39/NET4714 0 0.176433f
c_222 XI39/NET4774 0 0.176433f
c_223 XI39/NET6818 0 0.176433f
c_224 XI39/NET6690 0 0.176433f
c_225 XI39/NET8934 0 0.18066f
c_226 XI39/NET8994 0 0.176433f
c_227 XI39/NET8742 0 0.176433f
c_228 XI39/NET8682 0 0.176433f
c_229 XI39/NET9250 0 0.176433f
c_230 XI39/NET9190 0 0.176433f
c_231 XI39/NET9446 0 0.176433f
c_232 XI39/NET9506 0 0.176433f
c_233 XI39/NET8230 0 0.18066f
c_234 XI39/NET8170 0 0.176433f
c_235 XI39/NET8426 0 0.176433f
c_236 XI39/NET8486 0 0.176433f
c_237 XI39/NET7914 0 0.176433f
c_238 XI39/NET7974 0 0.176433f
c_239 XI39/NET7718 0 0.176433f
c_240 XI39/NET7658 0 0.176433f
c_241 XI39/NET10658 0 0.18066f
c_242 XI39/NET11222 0 0.176433f
c_243 XI39/NET10830 0 0.176433f
c_244 XI39/NET10890 0 0.176433f
c_245 XI39/NET11534 0 0.176433f
c_246 XI39/NET11026 0 0.176433f
c_247 XI39/NET11346 0 0.176433f
c_248 XI39/NET11310 0 0.176433f
c_249 XI39/NET10470 0 0.18066f
c_250 XI39/NET10530 0 0.176433f
c_251 XI39/NET10282 0 0.176433f
c_252 XI39/NET10222 0 0.176433f
c_253 XI39/NET9782 0 0.176433f
c_254 XI39/NET9706 0 0.176433f
c_255 XI39/NET9958 0 0.176433f
c_256 XI39/NET10018 0 0.176433f
c_257 XI39/NET5642 0 0.176433f
c_258 XI39/NET5458 0 0.176433f
c_259 XI39/NET5710 0 0.176433f
c_260 XI39/NET3558 0 0.176433f
c_261 XI39/NET5202 0 0.176433f
c_262 XI39/NET5390 0 0.176433f
c_263 XI39/NET5134 0 0.176433f
c_264 XI39/NET4946 0 0.176433f
c_265 XI39/NET3922 0 0.176433f
c_266 XI39/NET4110 0 0.176433f
c_267 XI39/NET3854 0 0.176433f
c_268 XI39/NET3666 0 0.176433f
c_269 XI39/NET4366 0 0.176433f
c_270 XI39/NET4178 0 0.176433f
c_271 XI39/NET4434 0 0.176433f
c_272 XI39/NET4622 0 0.176433f
c_273 XI39/NET6118 0 0.176433f
c_274 XI39/NET7454 0 0.176433f
c_275 XI39/NET6050 0 0.176433f
c_276 XI39/NET5862 0 0.176433f
c_277 XI39/NET7134 0 0.176433f
c_278 XI39/NET7522 0 0.176433f
c_279 XI39/NET7202 0 0.176433f
c_280 XI39/NET7014 0 0.176433f
c_281 XI39/NET6410 0 0.176433f
c_282 XI39/NET6222 0 0.176433f
c_283 XI39/NET6478 0 0.176433f
c_284 XI39/NET6666 0 0.176433f
c_285 XI39/NET4690 0 0.176433f
c_286 XI39/NET4878 0 0.176433f
c_287 XI39/NET6922 0 0.176433f
c_288 XI39/NET6762 0 0.176433f
c_289 XI39/NET8914 0 0.176433f
c_290 XI39/NET9098 0 0.176433f
c_291 XI39/NET8846 0 0.176433f
c_292 XI39/NET8658 0 0.176433f
c_293 XI39/NET9354 0 0.176433f
c_294 XI39/NET9166 0 0.176433f
c_295 XI39/NET9422 0 0.176433f
c_296 XI39/NET9610 0 0.176433f
c_297 XI39/NET8334 0 0.176433f
c_298 XI39/NET8146 0 0.176433f
c_299 XI39/NET8402 0 0.176433f
c_300 XI39/NET8590 0 0.176433f
c_301 XI39/NET7890 0 0.176433f
c_302 XI39/NET8078 0 0.176433f
c_303 XI39/NET7822 0 0.176433f
c_304 XI39/NET7634 0 0.176433f
c_305 XI39/NET10738 0 0.176433f
c_306 XI39/NET11198 0 0.176433f
c_307 XI39/NET10806 0 0.176433f
c_308 XI39/NET10994 0 0.176433f
c_309 XI39/NET11518 0 0.176433f
c_310 XI39/NET11130 0 0.176433f
c_311 XI39/NET11450 0 0.176433f
c_312 XI39/NET11638 0 0.176433f
c_313 XI39/NET10450 0 0.176433f
c_314 XI39/NET10630 0 0.176433f
c_315 XI39/NET10382 0 0.176433f
c_316 XI39/NET10202 0 0.176433f
c_317 XI39/NET9866 0 0.176433f
c_318 XI39/NET9686 0 0.176433f
c_319 XI39/NET9938 0 0.176433f
c_320 XI39/NET10090 0 0.176434f
c_321 XI39/NET5582 0 0.180473f
c_322 XI39/NET5522 0 0.176433f
c_323 XI39/NET5774 0 0.176433f
c_324 XI39/NET3534 0 0.176433f
c_325 XI39/NET5266 0 0.176433f
c_326 XI39/NET5326 0 0.176433f
c_327 XI39/NET5070 0 0.176433f
c_328 XI39/NET5010 0 0.176433f
c_329 XI39/NET3986 0 0.18066f
c_330 XI39/NET4046 0 0.176433f
c_331 XI39/NET3790 0 0.176433f
c_332 XI39/NET3730 0 0.176433f
c_333 XI39/NET4302 0 0.176433f
c_334 XI39/NET4242 0 0.176433f
c_335 XI39/NET4498 0 0.176433f
c_336 XI39/NET4558 0 0.176433f
c_337 XI39/NET7330 0 0.18066f
c_338 XI39/NET7390 0 0.176433f
c_339 XI39/NET5986 0 0.176433f
c_340 XI39/NET5926 0 0.176433f
c_341 XI39/NET7070 0 0.176433f
c_342 XI39/NET7570 0 0.176433f
c_343 XI39/NET7266 0 0.176433f
c_344 XI39/NET7302 0 0.176433f
c_345 XI39/NET6346 0 0.18066f
c_346 XI39/NET6286 0 0.176433f
c_347 XI39/NET6542 0 0.176433f
c_348 XI39/NET6602 0 0.176433f
c_349 XI39/NET4754 0 0.176433f
c_350 XI39/NET4814 0 0.176433f
c_351 XI39/NET6858 0 0.176433f
c_352 XI39/NET6794 0 0.176433f
c_353 XI39/NET8974 0 0.18066f
c_354 XI39/NET9034 0 0.176433f
c_355 XI39/NET8782 0 0.176433f
c_356 XI39/NET8722 0 0.176433f
c_357 XI39/NET9290 0 0.176433f
c_358 XI39/NET9230 0 0.176433f
c_359 XI39/NET9486 0 0.176433f
c_360 XI39/NET9546 0 0.176433f
c_361 XI39/NET8270 0 0.18066f
c_362 XI39/NET8210 0 0.176433f
c_363 XI39/NET8466 0 0.176433f
c_364 XI39/NET8526 0 0.176433f
c_365 XI39/NET7954 0 0.176433f
c_366 XI39/NET8014 0 0.176433f
c_367 XI39/NET7758 0 0.176433f
c_368 XI39/NET7698 0 0.176433f
c_369 XI39/NET11282 0 0.18066f
c_370 XI39/NET11262 0 0.176433f
c_371 XI39/NET10870 0 0.176433f
c_372 XI39/NET10930 0 0.176433f
c_373 XI39/NET11574 0 0.176433f
c_374 XI39/NET11066 0 0.176433f
c_375 XI39/NET11386 0 0.176433f
c_376 XI39/NET11662 0 0.176433f
c_377 XI39/NET10510 0 0.18066f
c_378 XI39/NET10570 0 0.176433f
c_379 XI39/NET10322 0 0.176433f
c_380 XI39/NET10262 0 0.176433f
c_381 XI39/NET9806 0 0.176433f
c_382 XI39/NET9746 0 0.176433f
c_383 XI39/NET9998 0 0.176433f
c_384 XI39/NET10122 0 0.176433f
c_385 XI39/NET5634 0 0.176433f
c_386 XI39/NET5450 0 0.176433f
c_387 XI39/NET5702 0 0.176433f
c_388 XI39/NET3582 0 0.176433f
c_389 XI39/NET5194 0 0.176433f
c_390 XI39/NET5382 0 0.176433f
c_391 XI39/NET5126 0 0.176433f
c_392 XI39/NET4938 0 0.176433f
c_393 XI39/NET3914 0 0.176433f
c_394 XI39/NET4102 0 0.176433f
c_395 XI39/NET3846 0 0.176433f
c_396 XI39/NET3658 0 0.176433f
c_397 XI39/NET4358 0 0.176433f
c_398 XI39/NET4170 0 0.176433f
c_399 XI39/NET4426 0 0.176433f
c_400 XI39/NET4614 0 0.176433f
c_401 XI39/NET6110 0 0.176433f
c_402 XI39/NET7446 0 0.176433f
c_403 XI39/NET6042 0 0.176433f
c_404 XI39/NET5854 0 0.176433f
c_405 XI39/NET7126 0 0.176433f
c_406 XI39/NET7514 0 0.176433f
c_407 XI39/NET7194 0 0.176433f
c_408 XI39/NET7006 0 0.176433f
c_409 XI39/NET6402 0 0.176433f
c_410 XI39/NET6214 0 0.176433f
c_411 XI39/NET6470 0 0.176433f
c_412 XI39/NET6658 0 0.176433f
c_413 XI39/NET4682 0 0.176433f
c_414 XI39/NET4870 0 0.176433f
c_415 XI39/NET6914 0 0.176433f
c_416 XI39/NET6754 0 0.176433f
c_417 XI39/NET8906 0 0.176433f
c_418 XI39/NET9090 0 0.176433f
c_419 XI39/NET8838 0 0.176433f
c_420 XI39/NET8650 0 0.176433f
c_421 XI39/NET9346 0 0.176433f
c_422 XI39/NET9158 0 0.176433f
c_423 XI39/NET9414 0 0.176433f
c_424 XI39/NET9602 0 0.176433f
c_425 XI39/NET8326 0 0.176433f
c_426 XI39/NET8138 0 0.176433f
c_427 XI39/NET8394 0 0.176433f
c_428 XI39/NET8582 0 0.176433f
c_429 XI39/NET7882 0 0.176433f
c_430 XI39/NET8070 0 0.176433f
c_431 XI39/NET7814 0 0.176433f
c_432 XI39/NET7626 0 0.176433f
c_433 XI39/NET10730 0 0.176433f
c_434 XI39/NET11190 0 0.176433f
c_435 XI39/NET10798 0 0.176433f
c_436 XI39/NET10986 0 0.176433f
c_437 XI39/NET11510 0 0.176433f
c_438 XI39/NET11122 0 0.176433f
c_439 XI39/NET11442 0 0.176433f
c_440 XI39/NET11630 0 0.176433f
c_441 XI39/NET10442 0 0.176433f
c_442 XI39/NET10622 0 0.176433f
c_443 XI39/NET10374 0 0.176433f
c_444 XI39/NET10194 0 0.176433f
c_445 XI39/NET9858 0 0.176433f
c_446 XI39/NET9678 0 0.176433f
c_447 XI39/NET9930 0 0.176433f
c_448 XI39/NET10058 0 0.176434f
c_449 XI39/NET5550 0 0.180473f
c_450 XI39/NET5498 0 0.176433f
c_451 XI39/NET5750 0 0.176433f
c_452 XI39/NET3510 0 0.176433f
c_453 XI39/NET5242 0 0.176433f
c_454 XI39/NET5302 0 0.176433f
c_455 XI39/NET5046 0 0.176433f
c_456 XI39/NET4986 0 0.176433f
c_457 XI39/NET3962 0 0.18066f
c_458 XI39/NET4022 0 0.176433f
c_459 XI39/NET3766 0 0.176433f
c_460 XI39/NET3706 0 0.176433f
c_461 XI39/NET4278 0 0.176433f
c_462 XI39/NET4218 0 0.176433f
c_463 XI39/NET4474 0 0.176433f
c_464 XI39/NET4534 0 0.176433f
c_465 XI39/NET6158 0 0.18066f
c_466 XI39/NET7366 0 0.176433f
c_467 XI39/NET5962 0 0.176433f
c_468 XI39/NET5902 0 0.176433f
c_469 XI39/NET7046 0 0.176433f
c_470 XI39/NET7546 0 0.176433f
c_471 XI39/NET7242 0 0.176433f
c_472 XI39/NET7278 0 0.176433f
c_473 XI39/NET6322 0 0.18066f
c_474 XI39/NET6262 0 0.176433f
c_475 XI39/NET6518 0 0.176433f
c_476 XI39/NET6578 0 0.176433f
c_477 XI39/NET4730 0 0.176433f
c_478 XI39/NET4790 0 0.176433f
c_479 XI39/NET6834 0 0.176433f
c_480 XI39/NET6706 0 0.176433f
c_481 XI39/NET8950 0 0.18066f
c_482 XI39/NET9010 0 0.176433f
c_483 XI39/NET8758 0 0.176433f
c_484 XI39/NET8698 0 0.176433f
c_485 XI39/NET9266 0 0.176433f
c_486 XI39/NET9206 0 0.176433f
c_487 XI39/NET9462 0 0.176433f
c_488 XI39/NET9522 0 0.176433f
c_489 XI39/NET8246 0 0.18066f
c_490 XI39/NET8186 0 0.176433f
c_491 XI39/NET8442 0 0.176433f
c_492 XI39/NET8502 0 0.176433f
c_493 XI39/NET7930 0 0.176433f
c_494 XI39/NET7990 0 0.176433f
c_495 XI39/NET7734 0 0.176433f
c_496 XI39/NET7674 0 0.176433f
c_497 XI39/NET10674 0 0.18066f
c_498 XI39/NET11238 0 0.176433f
c_499 XI39/NET10846 0 0.176433f
c_500 XI39/NET10906 0 0.176433f
c_501 XI39/NET11550 0 0.176433f
c_502 XI39/NET11042 0 0.176433f
c_503 XI39/NET11362 0 0.176433f
c_504 XI39/NET11326 0 0.176433f
c_505 XI39/NET10486 0 0.18066f
c_506 XI39/NET10546 0 0.176433f
c_507 XI39/NET10298 0 0.176433f
c_508 XI39/NET10238 0 0.176433f
c_509 XI39/NET9774 0 0.176433f
c_510 XI39/NET9722 0 0.176433f
c_511 XI39/NET9974 0 0.176433f
c_512 XI39/NET10034 0 0.176433f
c_513 XI39/NET5626 0 0.176433f
c_514 XI39/NET5442 0 0.176433f
c_515 XI39/NET5694 0 0.176433f
c_516 XI39/NET3550 0 0.176433f
c_517 XI39/NET5186 0 0.176433f
c_518 XI39/NET5374 0 0.176433f
c_519 XI39/NET5118 0 0.176433f
c_520 XI39/NET4930 0 0.176433f
c_521 XI39/NET3906 0 0.176433f
c_522 XI39/NET4094 0 0.176433f
c_523 XI39/NET3838 0 0.176433f
c_524 XI39/NET3650 0 0.176433f
c_525 XI39/NET4350 0 0.176433f
c_526 XI39/NET4162 0 0.176433f
c_527 XI39/NET4418 0 0.176433f
c_528 XI39/NET4606 0 0.176433f
c_529 XI39/NET6102 0 0.176433f
c_530 XI39/NET7438 0 0.176433f
c_531 XI39/NET6034 0 0.176433f
c_532 XI39/NET5846 0 0.176433f
c_533 XI39/NET7118 0 0.176433f
c_534 XI39/NET7506 0 0.176433f
c_535 XI39/NET7186 0 0.176433f
c_536 XI39/NET6998 0 0.176433f
c_537 XI39/NET6394 0 0.176433f
c_538 XI39/NET6206 0 0.176433f
c_539 XI39/NET6462 0 0.176433f
c_540 XI39/NET6650 0 0.176433f
c_541 XI39/NET4674 0 0.176433f
c_542 XI39/NET4862 0 0.176433f
c_543 XI39/NET6906 0 0.176433f
c_544 XI39/NET6746 0 0.176433f
c_545 XI39/NET8898 0 0.176433f
c_546 XI39/NET9082 0 0.176433f
c_547 XI39/NET8830 0 0.176433f
c_548 XI39/NET8642 0 0.176433f
c_549 XI39/NET9338 0 0.176433f
c_550 XI39/NET9150 0 0.176433f
c_551 XI39/NET9406 0 0.176433f
c_552 XI39/NET9594 0 0.176433f
c_553 XI39/NET8318 0 0.176433f
c_554 XI39/NET8130 0 0.176433f
c_555 XI39/NET8386 0 0.176433f
c_556 XI39/NET8574 0 0.176433f
c_557 XI39/NET7874 0 0.176433f
c_558 XI39/NET8062 0 0.176433f
c_559 XI39/NET7806 0 0.176433f
c_560 XI39/NET7618 0 0.176433f
c_561 XI39/NET10722 0 0.176433f
c_562 XI39/NET11182 0 0.176433f
c_563 XI39/NET10790 0 0.176433f
c_564 XI39/NET10978 0 0.176433f
c_565 XI39/NET11502 0 0.176433f
c_566 XI39/NET11114 0 0.176433f
c_567 XI39/NET11434 0 0.176433f
c_568 XI39/NET11622 0 0.176433f
c_569 XI39/NET10434 0 0.176433f
c_570 XI39/NET10614 0 0.176433f
c_571 XI39/NET10366 0 0.176433f
c_572 XI39/NET10186 0 0.176433f
c_573 XI39/NET9850 0 0.176433f
c_574 XI39/NET9670 0 0.176433f
c_575 XI39/NET9922 0 0.176433f
c_576 XI39/NET10082 0 0.176434f
c_577 XI39/NET5574 0 0.180473f
c_578 XI39/NET5490 0 0.176433f
c_579 XI39/NET5742 0 0.176433f
c_580 XI39/NET3502 0 0.176433f
c_581 XI39/NET5234 0 0.176433f
c_582 XI39/NET5294 0 0.176433f
c_583 XI39/NET5038 0 0.176433f
c_584 XI39/NET4978 0 0.176433f
c_585 XI39/NET3954 0 0.18066f
c_586 XI39/NET4014 0 0.176433f
c_587 XI39/NET3758 0 0.176433f
c_588 XI39/NET3698 0 0.176433f
c_589 XI39/NET4270 0 0.176433f
c_590 XI39/NET4210 0 0.176433f
c_591 XI39/NET4466 0 0.176433f
c_592 XI39/NET4526 0 0.176433f
c_593 XI39/NET6150 0 0.18066f
c_594 XI39/NET7358 0 0.176433f
c_595 XI39/NET5954 0 0.176433f
c_596 XI39/NET5894 0 0.176433f
c_597 XI39/NET7038 0 0.176433f
c_598 XI39/NET7538 0 0.176433f
c_599 XI39/NET7234 0 0.176433f
c_600 XI39/NET6958 0 0.176433f
c_601 XI39/NET6314 0 0.18066f
c_602 XI39/NET6254 0 0.176433f
c_603 XI39/NET6510 0 0.176433f
c_604 XI39/NET6570 0 0.176433f
c_605 XI39/NET4722 0 0.176433f
c_606 XI39/NET4782 0 0.176433f
c_607 XI39/NET6826 0 0.176433f
c_608 XI39/NET6698 0 0.176433f
c_609 XI39/NET8942 0 0.18066f
c_610 XI39/NET9002 0 0.176433f
c_611 XI39/NET8750 0 0.176433f
c_612 XI39/NET8690 0 0.176433f
c_613 XI39/NET9258 0 0.176433f
c_614 XI39/NET9198 0 0.176433f
c_615 XI39/NET9454 0 0.176433f
c_616 XI39/NET9514 0 0.176433f
c_617 XI39/NET8238 0 0.18066f
c_618 XI39/NET8178 0 0.176433f
c_619 XI39/NET8434 0 0.176433f
c_620 XI39/NET8494 0 0.176433f
c_621 XI39/NET7922 0 0.176433f
c_622 XI39/NET7982 0 0.176433f
c_623 XI39/NET7726 0 0.176433f
c_624 XI39/NET7666 0 0.176433f
c_625 XI39/NET10666 0 0.18066f
c_626 XI39/NET11230 0 0.176433f
c_627 XI39/NET10838 0 0.176433f
c_628 XI39/NET10898 0 0.176433f
c_629 XI39/NET11542 0 0.176433f
c_630 XI39/NET11034 0 0.176433f
c_631 XI39/NET11354 0 0.176433f
c_632 XI39/NET11318 0 0.176433f
c_633 XI39/NET10478 0 0.18066f
c_634 XI39/NET10538 0 0.176433f
c_635 XI39/NET10290 0 0.176433f
c_636 XI39/NET10230 0 0.176433f
c_637 XI39/NET9798 0 0.176433f
c_638 XI39/NET9714 0 0.176433f
c_639 XI39/NET9966 0 0.176433f
c_640 XI39/NET10026 0 0.176433f
c_641 XI39/NET5618 0 0.176433f
c_642 XI39/NET5434 0 0.176433f
c_643 XI39/NET5686 0 0.176433f
c_644 XI39/NET3590 0 0.176433f
c_645 XI39/NET5178 0 0.176433f
c_646 XI39/NET5366 0 0.176433f
c_647 XI39/NET5110 0 0.176433f
c_648 XI39/NET4922 0 0.176433f
c_649 XI39/NET3898 0 0.176433f
c_650 XI39/NET4086 0 0.176433f
c_651 XI39/NET3830 0 0.176433f
c_652 XI39/NET3642 0 0.176433f
c_653 XI39/NET4342 0 0.176433f
c_654 XI39/NET4154 0 0.176433f
c_655 XI39/NET4410 0 0.176433f
c_656 XI39/NET4598 0 0.176433f
c_657 XI39/NET6094 0 0.176433f
c_658 XI39/NET7430 0 0.176433f
c_659 XI39/NET6026 0 0.176433f
c_660 XI39/NET5838 0 0.176433f
c_661 XI39/NET7110 0 0.176433f
c_662 XI39/NET7498 0 0.176433f
c_663 XI39/NET7178 0 0.176433f
c_664 XI39/NET6990 0 0.176433f
c_665 XI39/NET6386 0 0.176433f
c_666 XI39/NET6198 0 0.176433f
c_667 XI39/NET6454 0 0.176433f
c_668 XI39/NET6642 0 0.176433f
c_669 XI39/NET4666 0 0.176433f
c_670 XI39/NET4854 0 0.176433f
c_671 XI39/NET6898 0 0.176433f
c_672 XI39/NET6738 0 0.176433f
c_673 XI39/NET8890 0 0.176433f
c_674 XI39/NET9074 0 0.176433f
c_675 XI39/NET8822 0 0.176433f
c_676 XI39/NET8634 0 0.176433f
c_677 XI39/NET9330 0 0.176433f
c_678 XI39/NET9142 0 0.176433f
c_679 XI39/NET9398 0 0.176433f
c_680 XI39/NET9586 0 0.176433f
c_681 XI39/NET8310 0 0.176433f
c_682 XI39/NET8122 0 0.176433f
c_683 XI39/NET8378 0 0.176433f
c_684 XI39/NET8566 0 0.176433f
c_685 XI39/NET7866 0 0.176433f
c_686 XI39/NET8054 0 0.176433f
c_687 XI39/NET7798 0 0.176433f
c_688 XI39/NET7610 0 0.176433f
c_689 XI39/NET10714 0 0.176433f
c_690 XI39/NET11174 0 0.176433f
c_691 XI39/NET10782 0 0.176433f
c_692 XI39/NET10970 0 0.176433f
c_693 XI39/NET11494 0 0.176433f
c_694 XI39/NET11106 0 0.176433f
c_695 XI39/NET11426 0 0.176433f
c_696 XI39/NET11614 0 0.176433f
c_697 XI39/NET10426 0 0.176433f
c_698 XI39/NET10606 0 0.176433f
c_699 XI39/NET10358 0 0.176433f
c_700 XI39/NET10178 0 0.176433f
c_701 XI39/NET9842 0 0.176433f
c_702 XI39/NET9662 0 0.176433f
c_703 XI39/NET9914 0 0.176433f
c_704 XI39/NET10050 0 0.176434f
c_705 XI39/NET5542 0 0.180473f
c_706 XI39/NET5514 0 0.176433f
c_707 XI39/NET5766 0 0.176433f
c_708 XI39/NET3526 0 0.176433f
c_709 XI39/NET5258 0 0.176433f
c_710 XI39/NET5318 0 0.176433f
c_711 XI39/NET5062 0 0.176433f
c_712 XI39/NET5002 0 0.176433f
c_713 XI39/NET3978 0 0.18066f
c_714 XI39/NET4038 0 0.176433f
c_715 XI39/NET3782 0 0.176433f
c_716 XI39/NET3722 0 0.176433f
c_717 XI39/NET4294 0 0.176433f
c_718 XI39/NET4234 0 0.176433f
c_719 XI39/NET4490 0 0.176433f
c_720 XI39/NET4550 0 0.176433f
c_721 XI39/NET7322 0 0.18066f
c_722 XI39/NET7382 0 0.176433f
c_723 XI39/NET5978 0 0.176433f
c_724 XI39/NET5918 0 0.176433f
c_725 XI39/NET7062 0 0.176433f
c_726 XI39/NET7562 0 0.176433f
c_727 XI39/NET7258 0 0.176433f
c_728 XI39/NET7294 0 0.176433f
c_729 XI39/NET6338 0 0.18066f
c_730 XI39/NET6278 0 0.176433f
c_731 XI39/NET6534 0 0.176433f
c_732 XI39/NET6594 0 0.176433f
c_733 XI39/NET4746 0 0.176433f
c_734 XI39/NET4806 0 0.176433f
c_735 XI39/NET6850 0 0.176433f
c_736 XI39/NET6786 0 0.176433f
c_737 XI39/NET8966 0 0.18066f
c_738 XI39/NET9026 0 0.176433f
c_739 XI39/NET8774 0 0.176433f
c_740 XI39/NET8714 0 0.176433f
c_741 XI39/NET9282 0 0.176433f
c_742 XI39/NET9222 0 0.176433f
c_743 XI39/NET9478 0 0.176433f
c_744 XI39/NET9538 0 0.176433f
c_745 XI39/NET8262 0 0.18066f
c_746 XI39/NET8202 0 0.176433f
c_747 XI39/NET8458 0 0.176433f
c_748 XI39/NET8518 0 0.176433f
c_749 XI39/NET7946 0 0.176433f
c_750 XI39/NET8006 0 0.176433f
c_751 XI39/NET7750 0 0.176433f
c_752 XI39/NET7690 0 0.176433f
c_753 XI39/NET11274 0 0.18066f
c_754 XI39/NET11254 0 0.176433f
c_755 XI39/NET10862 0 0.176433f
c_756 XI39/NET10922 0 0.176433f
c_757 XI39/NET11566 0 0.176433f
c_758 XI39/NET11058 0 0.176433f
c_759 XI39/NET11378 0 0.176433f
c_760 XI39/NET11654 0 0.176433f
c_761 XI39/NET10502 0 0.18066f
c_762 XI39/NET10562 0 0.176433f
c_763 XI39/NET10314 0 0.176433f
c_764 XI39/NET10254 0 0.176433f
c_765 XI39/NET9766 0 0.176433f
c_766 XI39/NET9738 0 0.176433f
c_767 XI39/NET9990 0 0.176433f
c_768 XI39/NET10114 0 0.176433f
c_769 XI39/NET5610 0 0.176433f
c_770 XI39/NET5426 0 0.176433f
c_771 XI39/NET5678 0 0.176433f
c_772 XI39/NET3598 0 0.176433f
c_773 XI39/NET5170 0 0.176433f
c_774 XI39/NET5358 0 0.176433f
c_775 XI39/NET5102 0 0.176433f
c_776 XI39/NET4914 0 0.176433f
c_777 XI39/NET3890 0 0.176433f
c_778 XI39/NET4078 0 0.176433f
c_779 XI39/NET3822 0 0.176433f
c_780 XI39/NET3634 0 0.176433f
c_781 XI39/NET4334 0 0.176433f
c_782 XI39/NET4146 0 0.176433f
c_783 XI39/NET4402 0 0.176433f
c_784 XI39/NET4590 0 0.176433f
c_785 XI39/NET6086 0 0.176433f
c_786 XI39/NET7422 0 0.176433f
c_787 XI39/NET6018 0 0.176433f
c_788 XI39/NET5830 0 0.176433f
c_789 XI39/NET7102 0 0.176433f
c_790 XI39/NET7490 0 0.176433f
c_791 XI39/NET7170 0 0.176433f
c_792 XI39/NET6982 0 0.176433f
c_793 XI39/NET6378 0 0.176433f
c_794 XI39/NET6190 0 0.176433f
c_795 XI39/NET6446 0 0.176433f
c_796 XI39/NET6634 0 0.176433f
c_797 XI39/NET4658 0 0.176433f
c_798 XI39/NET4846 0 0.176433f
c_799 XI39/NET6890 0 0.176433f
c_800 XI39/NET6730 0 0.176433f
c_801 XI39/NET8882 0 0.176433f
c_802 XI39/NET9066 0 0.176433f
c_803 XI39/NET8814 0 0.176433f
c_804 XI39/NET8626 0 0.176433f
c_805 XI39/NET9322 0 0.176433f
c_806 XI39/NET9134 0 0.176433f
c_807 XI39/NET9390 0 0.176433f
c_808 XI39/NET9578 0 0.176433f
c_809 XI39/NET8302 0 0.176433f
c_810 XI39/NET8114 0 0.176433f
c_811 XI39/NET8370 0 0.176433f
c_812 XI39/NET8558 0 0.176433f
c_813 XI39/NET7858 0 0.176433f
c_814 XI39/NET8046 0 0.176433f
c_815 XI39/NET7790 0 0.176433f
c_816 XI39/NET7602 0 0.176433f
c_817 XI39/NET10706 0 0.176433f
c_818 XI39/NET11166 0 0.176433f
c_819 XI39/NET10774 0 0.176433f
c_820 XI39/NET10962 0 0.176433f
c_821 XI39/NET11486 0 0.176433f
c_822 XI39/NET11098 0 0.176433f
c_823 XI39/NET11418 0 0.176433f
c_824 XI39/NET11606 0 0.176433f
c_825 XI39/NET10418 0 0.176433f
c_826 XI39/NET10598 0 0.176433f
c_827 XI39/NET10350 0 0.176433f
c_828 XI39/NET10170 0 0.176433f
c_829 XI39/NET9834 0 0.176433f
c_830 XI39/NET9654 0 0.176433f
c_831 XI39/NET9906 0 0.176433f
c_832 XI39/NET10074 0 0.176434f
c_833 XI39/NET5566 0 0.180473f
c_834 XI39/NET5506 0 0.176433f
c_835 XI39/NET5758 0 0.176433f
c_836 XI39/NET3518 0 0.176433f
c_837 XI39/NET5250 0 0.176433f
c_838 XI39/NET5310 0 0.176433f
c_839 XI39/NET5054 0 0.176433f
c_840 XI39/NET4994 0 0.176433f
c_841 XI39/NET3970 0 0.18066f
c_842 XI39/NET4030 0 0.176433f
c_843 XI39/NET3774 0 0.176433f
c_844 XI39/NET3714 0 0.176433f
c_845 XI39/NET4286 0 0.176433f
c_846 XI39/NET4226 0 0.176433f
c_847 XI39/NET4482 0 0.176433f
c_848 XI39/NET4542 0 0.176433f
c_849 XI39/NET6166 0 0.18066f
c_850 XI39/NET7374 0 0.176433f
c_851 XI39/NET5970 0 0.176433f
c_852 XI39/NET5910 0 0.176433f
c_853 XI39/NET7054 0 0.176433f
c_854 XI39/NET7554 0 0.176433f
c_855 XI39/NET7250 0 0.176433f
c_856 XI39/NET7286 0 0.176433f
c_857 XI39/NET6330 0 0.18066f
c_858 XI39/NET6270 0 0.176433f
c_859 XI39/NET6526 0 0.176433f
c_860 XI39/NET6586 0 0.176433f
c_861 XI39/NET4738 0 0.176433f
c_862 XI39/NET4798 0 0.176433f
c_863 XI39/NET6842 0 0.176433f
c_864 XI39/NET6778 0 0.176433f
c_865 XI39/NET8958 0 0.18066f
c_866 XI39/NET9018 0 0.176433f
c_867 XI39/NET8766 0 0.176433f
c_868 XI39/NET8706 0 0.176433f
c_869 XI39/NET9274 0 0.176433f
c_870 XI39/NET9214 0 0.176433f
c_871 XI39/NET9470 0 0.176433f
c_872 XI39/NET9530 0 0.176433f
c_873 XI39/NET8254 0 0.18066f
c_874 XI39/NET8194 0 0.176433f
c_875 XI39/NET8450 0 0.176433f
c_876 XI39/NET8510 0 0.176433f
c_877 XI39/NET7938 0 0.176433f
c_878 XI39/NET7998 0 0.176433f
c_879 XI39/NET7742 0 0.176433f
c_880 XI39/NET7682 0 0.176433f
c_881 XI39/NET10682 0 0.18066f
c_882 XI39/NET11246 0 0.176433f
c_883 XI39/NET10854 0 0.176433f
c_884 XI39/NET10914 0 0.176433f
c_885 XI39/NET11558 0 0.176433f
c_886 XI39/NET11050 0 0.176433f
c_887 XI39/NET11370 0 0.176433f
c_888 XI39/NET11334 0 0.176433f
c_889 XI39/NET10494 0 0.18066f
c_890 XI39/NET10554 0 0.176433f
c_891 XI39/NET10306 0 0.176433f
c_892 XI39/NET10246 0 0.176433f
c_893 XI39/NET9790 0 0.176433f
c_894 XI39/NET9730 0 0.176433f
c_895 XI39/NET9982 0 0.176433f
c_896 XI39/NET10106 0 0.176433f
c_897 XI39/NET5602 0 0.176433f
c_898 XI39/NET5418 0 0.176433f
c_899 XI39/NET5670 0 0.176433f
c_900 XI39/NET3606 0 0.176433f
c_901 XI39/NET5162 0 0.176433f
c_902 XI39/NET5350 0 0.176433f
c_903 XI39/NET5094 0 0.176433f
c_904 XI39/NET4906 0 0.176433f
c_905 XI39/NET3882 0 0.176433f
c_906 XI39/NET4070 0 0.176433f
c_907 XI39/NET3814 0 0.176433f
c_908 XI39/NET3626 0 0.176433f
c_909 XI39/NET4326 0 0.176433f
c_910 XI39/NET4138 0 0.176433f
c_911 XI39/NET4394 0 0.176433f
c_912 XI39/NET4582 0 0.176433f
c_913 XI39/NET6078 0 0.176433f
c_914 XI39/NET7414 0 0.176433f
c_915 XI39/NET6010 0 0.176433f
c_916 XI39/NET5822 0 0.176433f
c_917 XI39/NET7094 0 0.176433f
c_918 XI39/NET7482 0 0.176433f
c_919 XI39/NET7162 0 0.176433f
c_920 XI39/NET6974 0 0.176433f
c_921 XI39/NET6370 0 0.176433f
c_922 XI39/NET6182 0 0.176433f
c_923 XI39/NET6438 0 0.176433f
c_924 XI39/NET6626 0 0.176433f
c_925 XI39/NET4650 0 0.176433f
c_926 XI39/NET4838 0 0.176433f
c_927 XI39/NET6882 0 0.176433f
c_928 XI39/NET6722 0 0.176433f
c_929 XI39/NET8874 0 0.176433f
c_930 XI39/NET9058 0 0.176433f
c_931 XI39/NET8806 0 0.176433f
c_932 XI39/NET8618 0 0.176433f
c_933 XI39/NET9314 0 0.176433f
c_934 XI39/NET9126 0 0.176433f
c_935 XI39/NET9382 0 0.176433f
c_936 XI39/NET9570 0 0.176433f
c_937 XI39/NET8294 0 0.176433f
c_938 XI39/NET8106 0 0.176433f
c_939 XI39/NET8362 0 0.176433f
c_940 XI39/NET8550 0 0.176433f
c_941 XI39/NET7850 0 0.176433f
c_942 XI39/NET8038 0 0.176433f
c_943 XI39/NET7782 0 0.176433f
c_944 XI39/NET7594 0 0.176433f
c_945 XI39/NET10698 0 0.176433f
c_946 XI39/NET11158 0 0.176433f
c_947 XI39/NET10766 0 0.176433f
c_948 XI39/NET10954 0 0.176433f
c_949 XI39/NET11478 0 0.176433f
c_950 XI39/NET11090 0 0.176433f
c_951 XI39/NET11410 0 0.176433f
c_952 XI39/NET11598 0 0.176433f
c_953 XI39/NET10410 0 0.176433f
c_954 XI39/NET10590 0 0.176433f
c_955 XI39/NET10342 0 0.176433f
c_956 XI39/NET10162 0 0.176433f
c_957 XI39/NET9826 0 0.176433f
c_958 XI39/NET9646 0 0.176433f
c_959 XI39/NET9898 0 0.176433f
c_960 XI39/NET10042 0 0.176434f
c_961 XI39/NET5534 0 0.137954f
c_962 XI39/NET5474 0 0.136314f
c_963 XI39/NET5726 0 0.136314f
c_964 XI39/NET3486 0 0.136314f
c_965 XI39/NET5218 0 0.136314f
c_966 XI39/NET5278 0 0.136314f
c_967 XI39/NET5022 0 0.136314f
c_968 XI39/NET4962 0 0.136314f
c_969 XI39/NET3938 0 0.138908f
c_970 XI39/NET3998 0 0.136314f
c_971 XI39/NET3742 0 0.136314f
c_972 XI39/NET3682 0 0.136314f
c_973 XI39/NET4254 0 0.136314f
c_974 XI39/NET4194 0 0.136314f
c_975 XI39/NET4450 0 0.136314f
c_976 XI39/NET4510 0 0.136314f
c_977 XI39/NET6134 0 0.138908f
c_978 XI39/NET7342 0 0.136314f
c_979 XI39/NET5938 0 0.136314f
c_980 XI39/NET5878 0 0.136314f
c_981 XI39/NET5802 0 0.136314f
c_982 XI39/NET5790 0 0.136314f
c_983 XI39/NET7218 0 0.136314f
c_984 XI39/NET6942 0 0.136314f
c_985 XI39/NET6298 0 0.138908f
c_986 XI39/NET6238 0 0.136314f
c_987 XI39/NET6494 0 0.136314f
c_988 XI39/NET6554 0 0.136314f
c_989 XI39/NET4706 0 0.136314f
c_990 XI39/NET4766 0 0.136314f
c_991 XI39/NET6810 0 0.136314f
c_992 XI39/NET6682 0 0.136314f
c_993 XI39/NET8926 0 0.138908f
c_994 XI39/NET8986 0 0.136314f
c_995 XI39/NET8734 0 0.136314f
c_996 XI39/NET8674 0 0.136314f
c_997 XI39/NET9242 0 0.136314f
c_998 XI39/NET9182 0 0.136314f
c_999 XI39/NET9438 0 0.136314f
c_1000 XI39/NET9498 0 0.136314f
c_1001 XI39/NET8222 0 0.138908f
c_1002 XI39/NET8162 0 0.136314f
c_1003 XI39/NET8418 0 0.136314f
c_1004 XI39/NET8478 0 0.136314f
c_1005 XI39/NET7906 0 0.136314f
c_1006 XI39/NET7966 0 0.136314f
c_1007 XI39/NET7710 0 0.136314f
c_1008 XI39/NET7650 0 0.136314f
c_1009 XI39/NET10650 0 0.138908f
c_1010 XI39/NET11214 0 0.136314f
c_1011 XI39/NET10822 0 0.136314f
c_1012 XI39/NET10882 0 0.136314f
c_1013 XI39/NET11014 0 0.136314f
c_1014 XI39/NET11018 0 0.136314f
c_1015 XI39/NET11338 0 0.136314f
c_1016 XI39/NET11302 0 0.136314f
c_1017 XI39/NET10462 0 0.138908f
c_1018 XI39/NET10522 0 0.136314f
c_1019 XI39/NET10274 0 0.136314f
c_1020 XI39/NET10214 0 0.136314f
c_1021 XI39/NET9758 0 0.136314f
c_1022 XI39/NET9698 0 0.136314f
c_1023 XI39/NET9950 0 0.136314f
c_1024 XI39/NET10010 0 0.136314f
*
.include "ROM_TEST6.pex.spi.ROM_TEST6.pxi"
*
.ends
*
*
